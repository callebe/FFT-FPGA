library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT0 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT0;

architecture Behavioral of ROMFFT0 is

    signal Counter : integer range 0 to 1023 := 0;
	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 1 
	constant ROM_tb : ROM := (
		0 => "111000010100001010000",
		1 => "111000010100001010000",
		2 => "111000010100001010000",
		3 => "011000000101111110011",
		4 => "011000000101111110011",
		5 => "011000000101111110011",
		6 => "011010100100001110100",
		7 => "011010100100001110100",
		8 => "011010100100001110100",
		9 => "001010111100001010101",
		10 => "001010111100001010101",
		11 => "001010111100001010101",
		12 => "011001111100001010110",
		13 => "011001111100001010110",
		14 => "011001111100001010110",
		15 => "011001011101001010000",
		16 => "011001011101001010000",
		17 => "011001011101001010000",
		18 => "011000001101100010011",
		19 => "011000001101100010011",
		20 => "011000001101100010011",
		21 => "001000111100011110011",
		22 => "001000111100011110011",
		23 => "001000111100011110011",
		24 => "011000101100100010101",
		25 => "011000101100100010101",
		26 => "011000101100100010101",
		27 => "011000101100111010001",
		28 => "011000101100111010001",
		29 => "011000101100111010001",
		30 => "111011010100001010011",
		31 => "111011010100001010011",
		32 => "111011010100001010011",
		33 => "011001011100001010100",
		34 => "011001011100001010100",
		35 => "011001011100001010100",
		36 => "011001100100001110001",
		37 => "011001100100001110001",
		38 => "011001100100001110001",
		39 => "011000000101011010101",
		40 => "011000000101011010101",
		41 => "011000000101011010101",
		42 => "011010100100001010100",
		43 => "011010100100001010100",
		44 => "011010100100001010100",
		45 => "011011100100001110011",
		46 => "011011100100001110011",
		47 => "011011100100001110011",
		48 => "011000101100100110010",
		49 => "011000101100100110010",
		50 => "011000101100100110010",
		51 => "001001111100001010111",
		52 => "001001111100001010111",
		53 => "001001111100001010111",
		54 => "011010100100001110100",
		55 => "011010100100001110100",
		56 => "011010100100001110100",
		57 => "011010100100001010101",
		58 => "011010100100001010101",
		59 => "011010100100001010101",
		60 => "011011000100001110011",
		61 => "011011000100001110011",
		62 => "011011000100001110011",
		63 => "011010000100001010010",
		64 => "011010000100001010010",
		65 => "011010000100001010010",
		66 => "011000001101100010011",
		67 => "011000001101100010011",
		68 => "011000001101100010011",
		69 => "001000100100111010001",
		70 => "001000100100111010001",
		71 => "001000100100111010001",
		72 => "011000101100100010101",
		73 => "011000101100100010101",
		74 => "011000101100100010101",
		75 => "001000000100101110110",
		76 => "001000000100101110110",
		77 => "001000000100101110110",
		78 => "011000001101100010011",
		79 => "011000001101100010011",
		80 => "011000001101100010011",
		81 => "011010000100001110010",
		82 => "011010000100001110010",
		83 => "011010000100001110010",
		84 => "001000111100111010000",
		85 => "001000111100111010000",
		86 => "001000111100111010000",
		87 => "011000000101011010101",
		88 => "011000000101011010101",
		89 => "011000000101011010101",
		90 => "011010100100001010100",
		91 => "011010100100001010100",
		92 => "011010100100001010100",
		93 => "011000000101111010011",
		94 => "011000000101111010011",
		95 => "011000000101111010011",
		96 => "111000010100001010000",
		97 => "111000010100001010000",
		98 => "111000010100001010000",
		99 => "011010100100001110100",
		100 => "011010100100001110100",
		101 => "011010100100001110100",
		102 => "011001111100001010110",
		103 => "011001111100001010110",
		104 => "011001111100001010110",
		105 => "011000001101100010011",
		106 => "011000001101100010011",
		107 => "011000001101100010011",
		108 => "011000101100100010101",
		109 => "011000101100100010101",
		110 => "011000101100100010101",
		111 => "111011010100001010011",
		112 => "111011010100001010011",
		113 => "111011010100001010011",
		114 => "011001100100001110001",
		115 => "011001100100001110001",
		116 => "011001100100001110001",
		117 => "011010100100001010100",
		118 => "011010100100001010100",
		119 => "011010100100001010100",
		120 => "011000101100100110010",
		121 => "011000101100100110010",
		122 => "011000101100100110010",
		123 => "011010100100001110100",
		124 => "011010100100001110100",
		125 => "011010100100001110100",
		126 => "011011000100001110011",
		127 => "011011000100001110011",
		128 => "011011000100001110011",
		129 => "011000001101100010011",
		130 => "011000001101100010011",
		131 => "011000001101100010011",
		132 => "011000101100100010101",
		133 => "011000101100100010101",
		134 => "011000101100100010101",
		135 => "011000001101100010011",
		136 => "011000001101100010011",
		137 => "011000001101100010011",
		138 => "001000111100111010000",
		139 => "001000111100111010000",
		140 => "001000111100111010000",
		141 => "011010100100001010100",
		142 => "011010100100001010100",
		143 => "011010100100001010100",
		144 => "111000010100001010000",
		145 => "111000010100001010000",
		146 => "111000010100001010000",
		147 => "011010100100001110100",
		148 => "011010100100001110100",
		149 => "011010100100001110100",
		150 => "011001111100001010110",
		151 => "011001111100001010110",
		152 => "011001111100001010110",
		153 => "011000001101100010011",
		154 => "011000001101100010011",
		155 => "011000001101100010011",
		156 => "011000101100100010101",
		157 => "011000101100100010101",
		158 => "011000101100100010101",
		159 => "111011010100001010011",
		160 => "111011010100001010011",
		161 => "111011010100001010011",
		162 => "011001100100001110001",
		163 => "011001100100001110001",
		164 => "011001100100001110001",
		165 => "011010100100001010100",
		166 => "011010100100001010100",
		167 => "011010100100001010100",
		168 => "011000101100100110010",
		169 => "011000101100100110010",
		170 => "011000101100100110010",
		171 => "011010100100001110100",
		172 => "011010100100001110100",
		173 => "011010100100001110100",
		174 => "011011000100001110011",
		175 => "011011000100001110011",
		176 => "011011000100001110011",
		177 => "011000001101100010011",
		178 => "011000001101100010011",
		179 => "011000001101100010011",
		180 => "011000101100100010101",
		181 => "011000101100100010101",
		182 => "011000101100100010101",
		183 => "011000001101100010011",
		184 => "011000001101100010011",
		185 => "011000001101100010011",
		186 => "001000111100111010000",
		187 => "001000111100111010000",
		188 => "001000111100111010000",
		189 => "011010100100001010100",
		190 => "011010100100001010100",
		191 => "011010100100001010100",
		192 => "111000010100001010000",
		193 => "111000010100001010000",
		194 => "111000010100001010000",
		195 => "011001111100001010110",
		196 => "011001111100001010110",
		197 => "011001111100001010110",
		198 => "011000101100100010101",
		199 => "011000101100100010101",
		200 => "011000101100100010101",
		201 => "011001100100001110001",
		202 => "011001100100001110001",
		203 => "011001100100001110001",
		204 => "011000101100100110010",
		205 => "011000101100100110010",
		206 => "011000101100100110010",
		207 => "011011000100001110011",
		208 => "011011000100001110011",
		209 => "011011000100001110011",
		210 => "011000101100100010101",
		211 => "011000101100100010101",
		212 => "011000101100100010101",
		213 => "001000111100111010000",
		214 => "001000111100111010000",
		215 => "001000111100111010000",
		216 => "111000010100001010000",
		217 => "111000010100001010000",
		218 => "111000010100001010000",
		219 => "011001111100001010110",
		220 => "011001111100001010110",
		221 => "011001111100001010110",
		222 => "011000101100100010101",
		223 => "011000101100100010101",
		224 => "011000101100100010101",
		225 => "011001100100001110001",
		226 => "011001100100001110001",
		227 => "011001100100001110001",
		228 => "011000101100100110010",
		229 => "011000101100100110010",
		230 => "011000101100100110010",
		231 => "011011000100001110011",
		232 => "011011000100001110011",
		233 => "011011000100001110011",
		234 => "011000101100100010101",
		235 => "011000101100100010101",
		236 => "011000101100100010101",
		237 => "001000111100111010000",
		238 => "001000111100111010000",
		239 => "001000111100111010000",
		240 => "111000010100001010000",
		241 => "111000010100001010000",
		242 => "111000010100001010000",
		243 => "011001111100001010110",
		244 => "011001111100001010110",
		245 => "011001111100001010110",
		246 => "011000101100100010101",
		247 => "011000101100100010101",
		248 => "011000101100100010101",
		249 => "011001100100001110001",
		250 => "011001100100001110001",
		251 => "011001100100001110001",
		252 => "011000101100100110010",
		253 => "011000101100100110010",
		254 => "011000101100100110010",
		255 => "011011000100001110011",
		256 => "011011000100001110011",
		257 => "011011000100001110011",
		258 => "011000101100100010101",
		259 => "011000101100100010101",
		260 => "011000101100100010101",
		261 => "001000111100111010000",
		262 => "001000111100111010000",
		263 => "001000111100111010000",
		264 => "111000010100001010000",
		265 => "111000010100001010000",
		266 => "111000010100001010000",
		267 => "011001111100001010110",
		268 => "011001111100001010110",
		269 => "011001111100001010110",
		270 => "011000101100100010101",
		271 => "011000101100100010101",
		272 => "011000101100100010101",
		273 => "011001100100001110001",
		274 => "011001100100001110001",
		275 => "011001100100001110001",
		276 => "011000101100100110010",
		277 => "011000101100100110010",
		278 => "011000101100100110010",
		279 => "011011000100001110011",
		280 => "011011000100001110011",
		281 => "011011000100001110011",
		282 => "011000101100100010101",
		283 => "011000101100100010101",
		284 => "011000101100100010101",
		285 => "001000111100111010000",
		286 => "001000111100111010000",
		287 => "001000111100111010000",
		288 => "111000010100001010000",
		289 => "111000010100001010000",
		290 => "111000010100001010000",
		291 => "011000101100100010101",
		292 => "011000101100100010101",
		293 => "011000101100100010101",
		294 => "011000101100100110010",
		295 => "011000101100100110010",
		296 => "011000101100100110010",
		297 => "011000101100100010101",
		298 => "011000101100100010101",
		299 => "011000101100100010101",
		300 => "111000010100001010000",
		301 => "111000010100001010000",
		302 => "111000010100001010000",
		303 => "011000101100100010101",
		304 => "011000101100100010101",
		305 => "011000101100100010101",
		306 => "011000101100100110010",
		307 => "011000101100100110010",
		308 => "011000101100100110010",
		309 => "011000101100100010101",
		310 => "011000101100100010101",
		311 => "011000101100100010101",
		312 => "111000010100001010000",
		313 => "111000010100001010000",
		314 => "111000010100001010000",
		315 => "011000101100100010101",
		316 => "011000101100100010101",
		317 => "011000101100100010101",
		318 => "011000101100100110010",
		319 => "011000101100100110010",
		320 => "011000101100100110010",
		321 => "011000101100100010101",
		322 => "011000101100100010101",
		323 => "011000101100100010101",
		324 => "111000010100001010000",
		325 => "111000010100001010000",
		326 => "111000010100001010000",
		327 => "011000101100100010101",
		328 => "011000101100100010101",
		329 => "011000101100100010101",
		330 => "011000101100100110010",
		331 => "011000101100100110010",
		332 => "011000101100100110010",
		333 => "011000101100100010101",
		334 => "011000101100100010101",
		335 => "011000101100100010101",
		336 => "111000010100001010000",
		337 => "111000010100001010000",
		338 => "111000010100001010000",
		339 => "011000101100100010101",
		340 => "011000101100100010101",
		341 => "011000101100100010101",
		342 => "011000101100100110010",
		343 => "011000101100100110010",
		344 => "011000101100100110010",
		345 => "011000101100100010101",
		346 => "011000101100100010101",
		347 => "011000101100100010101",
		348 => "111000010100001010000",
		349 => "111000010100001010000",
		350 => "111000010100001010000",
		351 => "011000101100100010101",
		352 => "011000101100100010101",
		353 => "011000101100100010101",
		354 => "011000101100100110010",
		355 => "011000101100100110010",
		356 => "011000101100100110010",
		357 => "011000101100100010101",
		358 => "011000101100100010101",
		359 => "011000101100100010101",
		360 => "111000010100001010000",
		361 => "111000010100001010000",
		362 => "111000010100001010000",
		363 => "011000101100100010101",
		364 => "011000101100100010101",
		365 => "011000101100100010101",
		366 => "011000101100100110010",
		367 => "011000101100100110010",
		368 => "011000101100100110010",
		369 => "011000101100100010101",
		370 => "011000101100100010101",
		371 => "011000101100100010101",
		372 => "111000010100001010000",
		373 => "111000010100001010000",
		374 => "111000010100001010000",
		375 => "011000101100100010101",
		376 => "011000101100100010101",
		377 => "011000101100100010101",
		378 => "011000101100100110010",
		379 => "011000101100100110010",
		380 => "011000101100100110010",
		381 => "011000101100100010101",
		382 => "011000101100100010101",
		383 => "011000101100100010101",
		384 => "111000010100001010000",
		385 => "111000010100001010000",
		386 => "111000010100001010000",
		387 => "011000101100100110010",
		388 => "011000101100100110010",
		389 => "011000101100100110010",
		390 => "111000010100001010000",
		391 => "111000010100001010000",
		392 => "111000010100001010000",
		393 => "011000101100100110010",
		394 => "011000101100100110010",
		395 => "011000101100100110010",
		396 => "111000010100001010000",
		397 => "111000010100001010000",
		398 => "111000010100001010000",
		399 => "011000101100100110010",
		400 => "011000101100100110010",
		401 => "011000101100100110010",
		402 => "111000010100001010000",
		403 => "111000010100001010000",
		404 => "111000010100001010000",
		405 => "011000101100100110010",
		406 => "011000101100100110010",
		407 => "011000101100100110010",
		408 => "111000010100001010000",
		409 => "111000010100001010000",
		410 => "111000010100001010000",
		411 => "011000101100100110010",
		412 => "011000101100100110010",
		413 => "011000101100100110010",
		414 => "111000010100001010000",
		415 => "111000010100001010000",
		416 => "111000010100001010000",
		417 => "011000101100100110010",
		418 => "011000101100100110010",
		419 => "011000101100100110010",
		420 => "111000010100001010000",
		421 => "111000010100001010000",
		422 => "111000010100001010000",
		423 => "011000101100100110010",
		424 => "011000101100100110010",
		425 => "011000101100100110010",
		426 => "111000010100001010000",
		427 => "111000010100001010000",
		428 => "111000010100001010000",
		429 => "011000101100100110010",
		430 => "011000101100100110010",
		431 => "011000101100100110010",
		432 => "111000010100001010000",
		433 => "111000010100001010000",
		434 => "111000010100001010000",
		435 => "011000101100100110010",
		436 => "011000101100100110010",
		437 => "011000101100100110010",
		438 => "111000010100001010000",
		439 => "111000010100001010000",
		440 => "111000010100001010000",
		441 => "011000101100100110010",
		442 => "011000101100100110010",
		443 => "011000101100100110010",
		444 => "111000010100001010000",
		445 => "111000010100001010000",
		446 => "111000010100001010000",
		447 => "011000101100100110010",
		448 => "011000101100100110010",
		449 => "011000101100100110010",
		450 => "111000010100001010000",
		451 => "111000010100001010000",
		452 => "111000010100001010000",
		453 => "011000101100100110010",
		454 => "011000101100100110010",
		455 => "011000101100100110010",
		456 => "111000010100001010000",
		457 => "111000010100001010000",
		458 => "111000010100001010000",
		459 => "011000101100100110010",
		460 => "011000101100100110010",
		461 => "011000101100100110010",
		462 => "111000010100001010000",
		463 => "111000010100001010000",
		464 => "111000010100001010000",
		465 => "011000101100100110010",
		466 => "011000101100100110010",
		467 => "011000101100100110010",
		468 => "111000010100001010000",
		469 => "111000010100001010000",
		470 => "111000010100001010000",
		471 => "011000101100100110010",
		472 => "011000101100100110010",
		473 => "011000101100100110010",
		474 => "111000010100001010000",
		475 => "111000010100001010000",
		476 => "111000010100001010000",
		477 => "011000101100100110010",
		478 => "011000101100100110010",
		479 => "011000101100100110010",
		480 => "111000010100001010000",
		481 => "111000010100001010000",
		482 => "111000010100001010000",
		483 => "111000010100001010000",
		484 => "111000010100001010000",
		485 => "111000010100001010000",
		486 => "111000010100001010000",
		487 => "111000010100001010000",
		488 => "111000010100001010000",
		489 => "111000010100001010000",
		490 => "111000010100001010000",
		491 => "111000010100001010000",
		492 => "111000010100001010000",
		493 => "111000010100001010000",
		494 => "111000010100001010000",
		495 => "111000010100001010000",
		496 => "111000010100001010000",
		497 => "111000010100001010000",
		498 => "111000010100001010000",
		499 => "111000010100001010000",
		500 => "111000010100001010000",
		501 => "111000010100001010000",
		502 => "111000010100001010000",
		503 => "111000010100001010000",
		504 => "111000010100001010000",
		505 => "111000010100001010000",
		506 => "111000010100001010000",
		507 => "111000010100001010000",
		508 => "111000010100001010000",
		509 => "111000010100001010000",
		510 => "111000010100001010000",
		511 => "111000010100001010000",
		512 => "111000010100001010000",
		513 => "111000010100001010000",
		514 => "111000010100001010000",
		515 => "111000010100001010000",
		516 => "111000010100001010000",
		517 => "111000010100001010000",
		518 => "111000010100001010000",
		519 => "111000010100001010000",
		520 => "111000010100001010000",
		521 => "111000010100001010000",
		522 => "111000010100001010000",
		523 => "111000010100001010000",
		524 => "111000010100001010000",
		525 => "111000010100001010000",
		526 => "111000010100001010000",
		527 => "111000010100001010000",
		528 => "111000010100001010000",
		529 => "111000010100001010000",
		530 => "111000010100001010000",
		531 => "111000010100001010000",
		532 => "111000010100001010000",
		533 => "111000010100001010000",
		534 => "111000010100001010000",
		535 => "111000010100001010000",
		536 => "111000010100001010000",
		537 => "111000010100001010000",
		538 => "111000010100001010000",
		539 => "111000010100001010000",
		540 => "111000010100001010000",
		541 => "111000010100001010000",
		542 => "111000010100001010000",
		543 => "111000010100001010000",
		544 => "111000010100001010000",
		545 => "111000010100001010000",
		546 => "111000010100001010000",
		547 => "111000010100001010000",
		548 => "111000010100001010000",
		549 => "111000010100001010000",
		550 => "111000010100001010000",
		551 => "111000010100001010000",
		552 => "111000010100001010000",
		553 => "111000010100001010000",
		554 => "111000010100001010000",
		555 => "111000010100001010000",
		556 => "111000010100001010000",
		557 => "111000010100001010000",
		558 => "111000010100001010000",
		559 => "111000010100001010000",
		560 => "111000010100001010000",
		561 => "111000010100001010000",
		562 => "111000010100001010000",
		563 => "111000010100001010000",
		564 => "111000010100001010000",
		565 => "111000010100001010000",
		566 => "111000010100001010000",
		567 => "111000010100001010000",
		568 => "111000010100001010000",
		569 => "111000010100001010000",
		570 => "111000010100001010000",
		571 => "111000010100001010000",
		572 => "111000010100001010000",
		573 => "111000010100001010000",
		574 => "111000010100001010000",
		575 => "111000010100001010000",
		576 => "111000010100001010000",
		577 => "111000010100001010000",
		578 => "111000010100001010000",
		579 => "111000010100001010000",
		580 => "111000010100001010000",
		581 => "111000010100001010000",
		582 => "111000010100001010000",
		583 => "111000010100001010000",
		584 => "111000010100001010000",
		585 => "111000010100001010000",
		586 => "111000010100001010000",
		587 => "111000010100001010000",
		588 => "111000010100001010000",
		589 => "111000010100001010000",
		590 => "111000010100001010000",
		591 => "111000010100001010000",
		592 => "111000010100001010000",
		593 => "111000010100001010000",
		594 => "111000010100001010000",
		595 => "111000010100001010000",
		596 => "111000010100001010000",
		597 => "111000010100001010000",
		598 => "111000010100001010000",
		599 => "111000010100001010000",
		600 => "111000010100001010000",
		601 => "111000010100001010000",
		602 => "111000010100001010000",
		603 => "111000010100001010000",
		604 => "111000010100001010000",
		605 => "111000010100001010000",
		606 => "111000010100001010000",
		607 => "111000010100001010000",
		608 => "111000010100001010000",
		609 => "111000010100001010000",
		610 => "111000010100001010000",
		611 => "111000010100001010000",
		612 => "111000010100001010000",
		613 => "111000010100001010000",
		614 => "111000010100001010000",
		615 => "111000010100001010000",
		616 => "111000010100001010000",
		617 => "111000010100001010000",
		618 => "111000010100001010000",
		619 => "111000010100001010000",
		620 => "111000010100001010000",
		621 => "111000010100001010000",
		622 => "111000010100001010000",
		623 => "111000010100001010000",
		624 => "111000010100001010000",
		625 => "111000010100001010000",
		626 => "111000010100001010000",
		627 => "111000010100001010000",
		628 => "111000010100001010000",
		629 => "111000010100001010000",
		630 => "111000010100001010000",
		631 => "111000010100001010000",
		632 => "111000010100001010000",
		633 => "111000010100001010000",
		634 => "111000010100001010000",
		635 => "111000010100001010000",
		636 => "111000010100001010000",
		637 => "111000010100001010000",
		638 => "111000010100001010000",
		639 => "111000010100001010000",
		640 => "111000010100001010000",
		641 => "111000010100001010000",
		642 => "111000010100001010000",
		643 => "111000010100001010000",
		644 => "111000010100001010000",
		645 => "111000010100001010000",
		646 => "111000010100001010000",
		647 => "111000010100001010000",
		648 => "111000010100001010000",
		649 => "111000010100001010000",
		650 => "111000010100001010000",
		651 => "111000010100001010000",
		652 => "111000010100001010000",
		653 => "111000010100001010000",
		654 => "111000010100001010000",
		655 => "111000010100001010000",
		656 => "111000010100001010000",
		657 => "111000010100001010000",
		658 => "111000010100001010000",
		659 => "111000010100001010000",
		660 => "111000010100001010000",
		661 => "111000010100001010000",
		662 => "111000010100001010000",
		663 => "111000010100001010000",
		664 => "111000010100001010000",
		665 => "111000010100001010000",
		666 => "111000010100001010000",
		667 => "111000010100001010000",
		668 => "111000010100001010000",
		669 => "111000010100001010000",
		670 => "111000010100001010000",
		671 => "111000010100001010000",
		672 => "111000010100001010000",
		673 => "111000010100001010000",
		674 => "111000010100001010000",
		675 => "111000010100001010000",
		676 => "111000010100001010000",
		677 => "111000010100001010000",
		678 => "111000010100001010000",
		679 => "111000010100001010000",
		680 => "111000010100001010000",
		681 => "111000010100001010000",
		682 => "111000010100001010000",
		683 => "111000010100001010000",
		684 => "111000010100001010000",
		685 => "111000010100001010000",
		686 => "111000010100001010000",
		687 => "111000010100001010000",
		688 => "111000010100001010000",
		689 => "111000010100001010000",
		690 => "111000010100001010000",
		691 => "111000010100001010000",
		692 => "111000010100001010000",
		693 => "111000010100001010000",
		694 => "111000010100001010000",
		695 => "111000010100001010000",
		696 => "111000010100001010000",
		697 => "111000010100001010000",
		698 => "111000010100001010000",
		699 => "111000010100001010000",
		700 => "111000010100001010000",
		701 => "111000010100001010000",
		702 => "111000010100001010000",
		703 => "111000010100001010000",
		704 => "111000010100001010000",
		705 => "111000010100001010000",
		706 => "111000010100001010000",
		707 => "111000010100001010000",
		708 => "111000010100001010000",
		709 => "111000010100001010000",
		710 => "111000010100001010000",
		711 => "111000010100001010000",
		712 => "111000010100001010000",
		713 => "111000010100001010000",
		714 => "111000010100001010000",
		715 => "111000010100001010000",
		716 => "111000010100001010000",
		717 => "111000010100001010000",
		718 => "111000010100001010000",
		719 => "111000010100001010000",
		720 => "111000010100001010000",
		721 => "111000010100001010000",
		722 => "111000010100001010000",
		723 => "111000010100001010000",
		724 => "111000010100001010000",
		725 => "111000010100001010000",
		726 => "111000010100001010000",
		727 => "111000010100001010000",
		728 => "111000010100001010000",
		729 => "111000010100001010000",
		730 => "111000010100001010000",
		731 => "111000010100001010000",
		732 => "111000010100001010000",
		733 => "111000010100001010000",
		734 => "111000010100001010000",
		735 => "111000010100001010000",
		736 => "111000010100001010000",
		737 => "111000010100001010000",
		738 => "111000010100001010000",
		739 => "111000010100001010000",
		740 => "111000010100001010000",
		741 => "111000010100001010000",
		742 => "111000010100001010000",
		743 => "111000010100001010000",
		744 => "111000010100001010000",
		745 => "111000010100001010000",
		746 => "111000010100001010000",
		747 => "111000010100001010000",
		748 => "111000010100001010000",
		749 => "111000010100001010000",
		750 => "111000010100001010000",
		751 => "111000010100001010000",
		752 => "111000010100001010000",
		753 => "111000010100001010000",
		754 => "111000010100001010000",
		755 => "111000010100001010000",
		756 => "111000010100001010000",
		757 => "111000010100001010000",
		758 => "111000010100001010000",
		759 => "111000010100001010000",
		760 => "111000010100001010000",
		761 => "111000010100001010000",
		762 => "111000010100001010000",
		763 => "111000010100001010000",
		764 => "111000010100001010000",
		765 => "111000010100001010000",
		766 => "111000010100001010000",
		767 => "111000010100001010000",
		768 => "111000010100001010000",
		769 => "111000010100001010000",
		770 => "111000010100001010000",
		771 => "111000010100001010000",
		772 => "111000010100001010000",
		773 => "111000010100001010000",
		774 => "111000010100001010000",
		775 => "111000010100001010000",
		776 => "111000010100001010000",
		777 => "111000010100001010000",
		778 => "111000010100001010000",
		779 => "111000010100001010000",
		780 => "111000010100001010000",
		781 => "111000010100001010000",
		782 => "111000010100001010000",
		783 => "111000010100001010000",
		784 => "111000010100001010000",
		785 => "111000010100001010000",
		786 => "111000010100001010000",
		787 => "111000010100001010000",
		788 => "111000010100001010000",
		789 => "111000010100001010000",
		790 => "111000010100001010000",
		791 => "111000010100001010000",
		792 => "111000010100001010000",
		793 => "111000010100001010000",
		794 => "111000010100001010000",
		795 => "111000010100001010000",
		796 => "111000010100001010000",
		797 => "111000010100001010000",
		798 => "111000010100001010000",
		799 => "111000010100001010000",
		800 => "111000010100001010000",
		801 => "111000010100001010000",
		802 => "111000010100001010000",
		803 => "111000010100001010000",
		804 => "111000010100001010000",
		805 => "111000010100001010000",
		806 => "111000010100001010000",
		807 => "111000010100001010000",
		808 => "111000010100001010000",
		809 => "111000010100001010000",
		810 => "111000010100001010000",
		811 => "111000010100001010000",
		812 => "111000010100001010000",
		813 => "111000010100001010000",
		814 => "111000010100001010000",
		815 => "111000010100001010000",
		816 => "111000010100001010000",
		817 => "111000010100001010000",
		818 => "111000010100001010000",
		819 => "111000010100001010000",
		820 => "111000010100001010000",
		821 => "111000010100001010000",
		822 => "111000010100001010000",
		823 => "111000010100001010000",
		824 => "111000010100001010000",
		825 => "111000010100001010000",
		826 => "111000010100001010000",
		827 => "111000010100001010000",
		828 => "111000010100001010000",
		829 => "111000010100001010000",
		830 => "111000010100001010000",
		831 => "111000010100001010000",
		832 => "111000010100001010000",
		833 => "111000010100001010000",
		834 => "111000010100001010000",
		835 => "111000010100001010000",
		836 => "111000010100001010000",
		837 => "111000010100001010000",
		838 => "111000010100001010000",
		839 => "111000010100001010000",
		840 => "111000010100001010000",
		841 => "111000010100001010000",
		842 => "111000010100001010000",
		843 => "111000010100001010000",
		844 => "111000010100001010000",
		845 => "111000010100001010000",
		846 => "111000010100001010000",
		847 => "111000010100001010000",
		848 => "111000010100001010000",
		849 => "111000010100001010000",
		850 => "111000010100001010000",
		851 => "111000010100001010000",
		852 => "111000010100001010000",
		853 => "111000010100001010000",
		854 => "111000010100001010000",
		855 => "111000010100001010000",
		856 => "111000010100001010000",
		857 => "111000010100001010000",
		858 => "111000010100001010000",
		859 => "111000010100001010000",
		860 => "111000010100001010000",
		861 => "111000010100001010000",
		862 => "111000010100001010000",
		863 => "111000010100001010000");

begin

    --Output
    Data <= Rom_tb(Counter);
    
    --Process to acess Data
    process(Adress, reset)
    
    begin
    
        if(reset = '1')then
            Counter <= 0;
        
        elsif(Adress'event and Adress = '1') then
            if(Counter < 863) then
                Counter <= Counter + 1;
            end if;
        
        end if;
    
    end process;

end Behavioral;