--------------------------------------------------------------------
--------------------------------------------------------------------
--                                                                --
--                       Recep��o UART                            --
--    O clock usado na recep��o est� a 153600 Hz, exatamente 16   --
-- vezes maior que a velocidade de transmiss�o (9600 Hz). Para    --
-- que assim possa notar as mudan�as no sinal durante o ciclo do  --   
-- sinal de 9600 Hz com resolu��o de 16 pontos.                   --
--                                                                --
--       clk -> 153600 Hz                                           --
--			ActiveTx -> Sinal que aciona a trasmiss�o                --
--       DataTx -> Informa��o � transmitir                        --
--       Tx -> Bit de transmiss�o serial                          --
--       FinishTx -> Sinal que marca o fim da trasmiss�o          --
--                                                                --
--------------------------------------------------------------------
--------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_unsigned.ALL;
USE IEEE.numeric_std.ALL;
USE work.MainPackage.ALL;

ENTITY UARTRx IS
	PORT(clk : IN STD_LOGIC;
		reset : IN STD_LOGIC;
		Rx : IN STD_LOGIC;
		DataRx : OUT STD_LOGIC_VECTOR(7 downto 0);
		FinishRx : OUT STD_LOGIC);
END UARTRx;

ARCHITECTURE Logic OF UARTRx IS

	TYPE State IS (ResetRx, IdleRx, SendRx, StopRx);
	SIGNAL CurrentState : State := IdleRx;
	SIGNAL NextState : State := IdleRx;
	SIGNAL CounterData : INTEGER  RANGE 7 DOWNTO 0 := 0;
	SIGNAL FilterRx : STD_LOGIC := '1';
	SIGNAL CurrentStateRx : INTEGER  RANGE 3 DOWNTO 0 := 3;
	TYPE TestTYPE IS ARRAY(15 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
	
BEGIN

	---------------------------------------------------------------
	--              Filtro do Sinal de Entrada Rx                --
	---------------------------------------------------------------
	FilterStateMachine : PROCESS(clk, reset)
	
	BEGIN
	
		IF(reset = '1') THEN
			FilterRx <= '1';
			CurrentStateRx <= 3;
		
		ELSIF(clk = '1' AND clk'event) THEN
			IF(Rx = '0' AND CurrentStateRx /= 0) THEN
				IF(CurrentStateRx = 1) THEN
					FilterRx <= '0';
				
				END IF;
				CurrentStateRx <= CurrentStateRx - 1;
			
			ELSIF(Rx = '1' AND CurrentStateRx /= 3) then
				IF(CurrentStateRx = 2) THEN
					FilterRx <= '1';
			
				END IF;
				CurrentStateRx <= CurrentStateRx + 1;
			
			END IF;
		
		END IF;
	
	END PROCESS;
	
	---------------------------------------------------------------
	--                   Atualiza��o de Estatos                  --
	---------------------------------------------------------------
	UpdateState : PROCESS(clk, reset)
	
		VARIABLE Ping : INTEGER RANGE 15 DOWNTO 0 := 0;
		VARIABLE DataRxBuffer : STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');

	BEGIN
	
		IF(reset = '1') THEN
			Ping := 0;
			CurrentState <= ResetRx;
			CounterData  <= 0;
			DataRxBuffer := "00000000";
		
		ELSIF(clk = '1' AND clk'event) THEN
			IF(Ping = 15 OR (CurrentState = IdleRx AND NextState = SendRx AND Ping = 7) OR (CurrentState = IdleRx AND NextState = IdleRx)) THEN
				Ping := 0;
				CurrentState <= NextState;
				IF(CurrentState = SendRx) THEN
					DataRxBuffer := Shifter(DataRxBuffer, 1,'0');
					DataRxBuffer(0)  :=  FilterRx;
					--DataRxBuffer = "01011010";
					CounterData <= CounterData + 1;
				
				ELSE
					DataRxBuffer := DataRxBuffer;
					CounterData <= 0;
					IF(CurrentState = StopRx) THEN
						DataRx <= DataRxBuffer;
						
					ELSIF(CurrentState = IdleRx) THEN
						DataRxBuffer := "00000000";
						
					END IF;
				END IF;
			
			ELSE
				DataRxBuffer := DataRxBuffer;
				CurrentState <= CurrentState;
				Ping := Ping + 1;
				
			END IF;
			
		END IF;
	 
	END PROCESS;

	---------------------------------------------------------------
	--                   M�quinas de Estados                     --
	---------------------------------------------------------------
	StateMachine : PROCESS(CurrentState, FilterRx, CounterData)
	
	BEGIN
	
		CASE CurrentState IS

			WHEN ResetRx =>
				FinishRx <= '0';
				NextState <= IdleRx;

			WHEN IdleRx =>
				FinishRx <= 'X';
				IF(FilterRx = '0') THEN
					NextState <= SendRx;
				
				ELSE
					NextState <= IdleRx;
				
				END IF;

			WHEN SendRx =>
				FinishRx <= '0';
				IF(CounterData = 7) THEN
					NextState <= StopRx;
				
				ELSE
					NextState <= SendRx;
				
				END IF;

			WHEN StopRx =>
				FinishRx <= '1';
				IF(FilterRx = '1') THEN
					NextState <= IdleRx;
				
				ELSE
					NextState <= StopRx;
				
				END IF;

			WHEN OTHERS =>
				FinishRx <= '0';
				NextState <= ResetRx;

		END CASE;
	  
	END PROCESS;
	 
END Logic;
