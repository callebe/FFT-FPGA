library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT7 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT7;

architecture Behavioral of ROMFFT7 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 8 
	constant ROM_tb : ROM := (
		0 => "001010100101111110000",
		1 => "001010100101111110000",
		2 => "001010100101111110000",
		3 => "011011100100001010110",
		4 => "011011100100001010110",
		5 => "011011100100001010110",
		6 => "011011111100001010101",
		7 => "011011111100001010101",
		8 => "011011111100001010101",
		9 => "011010100100101110000",
		10 => "011010100100101110000",
		11 => "011010100100101110000",
		12 => "011000110100001010101",
		13 => "011000110100001010101",
		14 => "011000110100001010101",
		15 => "011000111100111010000",
		16 => "011000111100111010000",
		17 => "011000111100111010000",
		18 => "011000000100111010000",
		19 => "011000000100111010000",
		20 => "011000000100111010000",
		21 => "011000101100111110001",
		22 => "011000101100111110001",
		23 => "011000101100111110001",
		24 => "001001011100111010000",
		25 => "001001011100111010000",
		26 => "001001011100111010000",
		27 => "011000111100011110011",
		28 => "011000111100011110011",
		29 => "011000111100011110011",
		30 => "011001111100001010100",
		31 => "011001111100001010100",
		32 => "011001111100001010100",
		33 => "011000001101100010011",
		34 => "011000001101100010011",
		35 => "011000001101100010011",
		36 => "011001000100001110001",
		37 => "011001000100001110001",
		38 => "011001000100001110001",
		39 => "011001011100001010101",
		40 => "011001011100001010101",
		41 => "011001011100001010101",
		42 => "011000000101101010011",
		43 => "011000000101101010011",
		44 => "011000000101101010011",
		45 => "011100100100001110100",
		46 => "011100100100001110100",
		47 => "011100100100001110100",
		48 => "011000000101010011010",
		49 => "011000000101010011010",
		50 => "011000000101010011010",
		51 => "011011100100001010110",
		52 => "011011100100001010110",
		53 => "011011100100001010110",
		54 => "011000001110010010101",
		55 => "011000001110010010101",
		56 => "011000001110010010101",
		57 => "001000011101011010010",
		58 => "001000011101011010010",
		59 => "001000011101011010010",
		60 => "001000111100001110101",
		61 => "001000111100001110101",
		62 => "001000111100001110101",
		63 => "011001100100001010001",
		64 => "011001100100001010001",
		65 => "011001100100001010001",
		66 => "011001100100001110000",
		67 => "011001100100001110000",
		68 => "011001100100001110000",
		69 => "001000111100011110011",
		70 => "001000111100011110011",
		71 => "001000111100011110011",
		72 => "001001011100111010000",
		73 => "001001011100111010000",
		74 => "001001011100111010000",
		75 => "001000100100111110001",
		76 => "001000100100111110001",
		77 => "001000100100111110001",
		78 => "011010000100001110011",
		79 => "011010000100001110011",
		80 => "011010000100001110011",
		81 => "011000001101100010011",
		82 => "011000001101100010011",
		83 => "011000001101100010011",
		84 => "001000111100101010000",
		85 => "001000111100101010000",
		86 => "001000111100101010000",
		87 => "011010100100001110010",
		88 => "011010100100001110010",
		89 => "011010100100001110010",
		90 => "011011000100001110011",
		91 => "011011000100001110011",
		92 => "011011000100001110011",
		93 => "001010011110011010000",
		94 => "001010011110011010000",
		95 => "001010011110011010000",
		96 => "011011100101001110000",
		97 => "011011100101001110000",
		98 => "011011100101001110000",
		99 => "001001111100001010101",
		100 => "001001111100001010101",
		101 => "001001111100001010101",
		102 => "001011011100001010011",
		103 => "001011011100001010011",
		104 => "001011011100001010011",
		105 => "001000111100011110011",
		106 => "001000111100011110011",
		107 => "001000111100011110011",
		108 => "011000001100101010101",
		109 => "011000001100101010101",
		110 => "011000001100101010101",
		111 => "011000000101011010010",
		112 => "011000000101011010010",
		113 => "011000000101011010010",
		114 => "011010100100001110100",
		115 => "011010100100001110100",
		116 => "011010100100001110100",
		117 => "011011011101111010000",
		118 => "011011011101111010000",
		119 => "011011011101111010000",
		120 => "001000011101111010100",
		121 => "001000011101111010100",
		122 => "001000011101111010100",
		123 => "011010100100001010011",
		124 => "011010100100001010011",
		125 => "011010100100001010011",
		126 => "011001100100001010110",
		127 => "011001100100001010110",
		128 => "011001100100001010110",
		129 => "001000100100111010001",
		130 => "001000100100111010001",
		131 => "001000100100111010001",
		132 => "001000100100111110001",
		133 => "001000100100111110001",
		134 => "001000100100111110001",
		135 => "011000000101011010010",
		136 => "011000000101011010010",
		137 => "011000000101011010010",
		138 => "011010100100001110100",
		139 => "011010100100001110100",
		140 => "011010100100001110100",
		141 => "011011100100001010110",
		142 => "011011100100001010110",
		143 => "011011100100001010110",
		144 => "011011100101001110000",
		145 => "011011100101001110000",
		146 => "011011100101001110000",
		147 => "001001111100001010101",
		148 => "001001111100001010101",
		149 => "001001111100001010101",
		150 => "001011011100001010011",
		151 => "001011011100001010011",
		152 => "001011011100001010011",
		153 => "001000111100011110011",
		154 => "001000111100011110011",
		155 => "001000111100011110011",
		156 => "011000001100101010101",
		157 => "011000001100101010101",
		158 => "011000001100101010101",
		159 => "011000000101011010010",
		160 => "011000000101011010010",
		161 => "011000000101011010010",
		162 => "011010100100001110100",
		163 => "011010100100001110100",
		164 => "011010100100001110100",
		165 => "011011011101111010000",
		166 => "011011011101111010000",
		167 => "011011011101111010000",
		168 => "001000011101111010100",
		169 => "001000011101111010100",
		170 => "001000011101111010100",
		171 => "011010100100001010011",
		172 => "011010100100001010011",
		173 => "011010100100001010011",
		174 => "011001100100001010110",
		175 => "011001100100001010110",
		176 => "011001100100001010110",
		177 => "001000100100111010001",
		178 => "001000100100111010001",
		179 => "001000100100111010001",
		180 => "001000100100111110001",
		181 => "001000100100111110001",
		182 => "001000100100111110001",
		183 => "011000000101011010010",
		184 => "011000000101011010010",
		185 => "011000000101011010010",
		186 => "011010100100001110100",
		187 => "011010100100001110100",
		188 => "011010100100001110100",
		189 => "011011100100001010110",
		190 => "011011100100001010110",
		191 => "011011100100001010110",
		192 => "001010011100001010111",
		193 => "001010011100001010111",
		194 => "001010011100001010111",
		195 => "001001011100001010100",
		196 => "001001011100001010100",
		197 => "001001011100001010100",
		198 => "001001111100011110010",
		199 => "001001111100011110010",
		200 => "001001111100011110010",
		201 => "011000000101011010010",
		202 => "011000000101011010010",
		203 => "011000000101011010010",
		204 => "001000011101101010011",
		205 => "001000011101101010011",
		206 => "001000011101101010011",
		207 => "011010000100001010010",
		208 => "011010000100001010010",
		209 => "011010000100001010010",
		210 => "011001000100001010011",
		211 => "011001000100001010011",
		212 => "011001000100001010011",
		213 => "001001011101011010000",
		214 => "001001011101011010000",
		215 => "001001011101011010000",
		216 => "001010011100001010111",
		217 => "001010011100001010111",
		218 => "001010011100001010111",
		219 => "001001011100001010100",
		220 => "001001011100001010100",
		221 => "001001011100001010100",
		222 => "001001111100011110010",
		223 => "001001111100011110010",
		224 => "001001111100011110010",
		225 => "011000000101011010010",
		226 => "011000000101011010010",
		227 => "011000000101011010010",
		228 => "001000011101101010011",
		229 => "001000011101101010011",
		230 => "001000011101101010011",
		231 => "011010000100001010010",
		232 => "011010000100001010010",
		233 => "011010000100001010010",
		234 => "011001000100001010011",
		235 => "011001000100001010011",
		236 => "011001000100001010011",
		237 => "001001011101011010000",
		238 => "001001011101011010000",
		239 => "001001011101011010000",
		240 => "001010011100001010111",
		241 => "001010011100001010111",
		242 => "001010011100001010111",
		243 => "001001011100001010100",
		244 => "001001011100001010100",
		245 => "001001011100001010100",
		246 => "001001111100011110010",
		247 => "001001111100011110010",
		248 => "001001111100011110010",
		249 => "011000000101011010010",
		250 => "011000000101011010010",
		251 => "011000000101011010010",
		252 => "001000011101101010011",
		253 => "001000011101101010011",
		254 => "001000011101101010011",
		255 => "011010000100001010010",
		256 => "011010000100001010010",
		257 => "011010000100001010010",
		258 => "011001000100001010011",
		259 => "011001000100001010011",
		260 => "011001000100001010011",
		261 => "001001011101011010000",
		262 => "001001011101011010000",
		263 => "001001011101011010000",
		264 => "001010011100001010111",
		265 => "001010011100001010111",
		266 => "001010011100001010111",
		267 => "001001011100001010100",
		268 => "001001011100001010100",
		269 => "001001011100001010100",
		270 => "001001111100011110010",
		271 => "001001111100011110010",
		272 => "001001111100011110010",
		273 => "011000000101011010010",
		274 => "011000000101011010010",
		275 => "011000000101011010010",
		276 => "001000011101101010011",
		277 => "001000011101101010011",
		278 => "001000011101101010011",
		279 => "011010000100001010010",
		280 => "011010000100001010010",
		281 => "011010000100001010010",
		282 => "011001000100001010011",
		283 => "011001000100001010011",
		284 => "011001000100001010011",
		285 => "001001011101011010000",
		286 => "001001011101011010000",
		287 => "001001011101011010000",
		288 => "001001111100001010101",
		289 => "001001111100001010101",
		290 => "001001111100001010101",
		291 => "011000001101110010011",
		292 => "011000001101110010011",
		293 => "011000001101110010011",
		294 => "001000011101011010010",
		295 => "001000011101011010010",
		296 => "001000011101011010010",
		297 => "011000001101110010011",
		298 => "011000001101110010011",
		299 => "011000001101110010011",
		300 => "001001111100001010101",
		301 => "001001111100001010101",
		302 => "001001111100001010101",
		303 => "011000001101110010011",
		304 => "011000001101110010011",
		305 => "011000001101110010011",
		306 => "001000011101011010010",
		307 => "001000011101011010010",
		308 => "001000011101011010010",
		309 => "011000001101110010011",
		310 => "011000001101110010011",
		311 => "011000001101110010011",
		312 => "001001111100001010101",
		313 => "001001111100001010101",
		314 => "001001111100001010101",
		315 => "011000001101110010011",
		316 => "011000001101110010011",
		317 => "011000001101110010011",
		318 => "001000011101011010010",
		319 => "001000011101011010010",
		320 => "001000011101011010010",
		321 => "011000001101110010011",
		322 => "011000001101110010011",
		323 => "011000001101110010011",
		324 => "001001111100001010101",
		325 => "001001111100001010101",
		326 => "001001111100001010101",
		327 => "011000001101110010011",
		328 => "011000001101110010011",
		329 => "011000001101110010011",
		330 => "001000011101011010010",
		331 => "001000011101011010010",
		332 => "001000011101011010010",
		333 => "011000001101110010011",
		334 => "011000001101110010011",
		335 => "011000001101110010011",
		336 => "001001111100001010101",
		337 => "001001111100001010101",
		338 => "001001111100001010101",
		339 => "011000001101110010011",
		340 => "011000001101110010011",
		341 => "011000001101110010011",
		342 => "001000011101011010010",
		343 => "001000011101011010010",
		344 => "001000011101011010010",
		345 => "011000001101110010011",
		346 => "011000001101110010011",
		347 => "011000001101110010011",
		348 => "001001111100001010101",
		349 => "001001111100001010101",
		350 => "001001111100001010101",
		351 => "011000001101110010011",
		352 => "011000001101110010011",
		353 => "011000001101110010011",
		354 => "001000011101011010010",
		355 => "001000011101011010010",
		356 => "001000011101011010010",
		357 => "011000001101110010011",
		358 => "011000001101110010011",
		359 => "011000001101110010011",
		360 => "001001111100001010101",
		361 => "001001111100001010101",
		362 => "001001111100001010101",
		363 => "011000001101110010011",
		364 => "011000001101110010011",
		365 => "011000001101110010011",
		366 => "001000011101011010010",
		367 => "001000011101011010010",
		368 => "001000011101011010010",
		369 => "011000001101110010011",
		370 => "011000001101110010011",
		371 => "011000001101110010011",
		372 => "001001111100001010101",
		373 => "001001111100001010101",
		374 => "001001111100001010101",
		375 => "011000001101110010011",
		376 => "011000001101110010011",
		377 => "011000001101110010011",
		378 => "001000011101011010010",
		379 => "001000011101011010010",
		380 => "001000011101011010010",
		381 => "011000001101110010011",
		382 => "011000001101110010011",
		383 => "011000001101110010011",
		384 => "001000111100011110011",
		385 => "001000111100011110011",
		386 => "001000111100011110011",
		387 => "001000100100111010001",
		388 => "001000100100111010001",
		389 => "001000100100111010001",
		390 => "001000111100011110011",
		391 => "001000111100011110011",
		392 => "001000111100011110011",
		393 => "001000100100111010001",
		394 => "001000100100111010001",
		395 => "001000100100111010001",
		396 => "001000111100011110011",
		397 => "001000111100011110011",
		398 => "001000111100011110011",
		399 => "001000100100111010001",
		400 => "001000100100111010001",
		401 => "001000100100111010001",
		402 => "001000111100011110011",
		403 => "001000111100011110011",
		404 => "001000111100011110011",
		405 => "001000100100111010001",
		406 => "001000100100111010001",
		407 => "001000100100111010001",
		408 => "001000111100011110011",
		409 => "001000111100011110011",
		410 => "001000111100011110011",
		411 => "001000100100111010001",
		412 => "001000100100111010001",
		413 => "001000100100111010001",
		414 => "001000111100011110011",
		415 => "001000111100011110011",
		416 => "001000111100011110011",
		417 => "001000100100111010001",
		418 => "001000100100111010001",
		419 => "001000100100111010001",
		420 => "001000111100011110011",
		421 => "001000111100011110011",
		422 => "001000111100011110011",
		423 => "001000100100111010001",
		424 => "001000100100111010001",
		425 => "001000100100111010001",
		426 => "001000111100011110011",
		427 => "001000111100011110011",
		428 => "001000111100011110011",
		429 => "001000100100111010001",
		430 => "001000100100111010001",
		431 => "001000100100111010001",
		432 => "001000111100011110011",
		433 => "001000111100011110011",
		434 => "001000111100011110011",
		435 => "001000100100111010001",
		436 => "001000100100111010001",
		437 => "001000100100111010001",
		438 => "001000111100011110011",
		439 => "001000111100011110011",
		440 => "001000111100011110011",
		441 => "001000100100111010001",
		442 => "001000100100111010001",
		443 => "001000100100111010001",
		444 => "001000111100011110011",
		445 => "001000111100011110011",
		446 => "001000111100011110011",
		447 => "001000100100111010001",
		448 => "001000100100111010001",
		449 => "001000100100111010001",
		450 => "001000111100011110011",
		451 => "001000111100011110011",
		452 => "001000111100011110011",
		453 => "001000100100111010001",
		454 => "001000100100111010001",
		455 => "001000100100111010001",
		456 => "001000111100011110011",
		457 => "001000111100011110011",
		458 => "001000111100011110011",
		459 => "001000100100111010001",
		460 => "001000100100111010001",
		461 => "001000100100111010001",
		462 => "001000111100011110011",
		463 => "001000111100011110011",
		464 => "001000111100011110011",
		465 => "001000100100111010001",
		466 => "001000100100111010001",
		467 => "001000100100111010001",
		468 => "001000111100011110011",
		469 => "001000111100011110011",
		470 => "001000111100011110011",
		471 => "001000100100111010001",
		472 => "001000100100111010001",
		473 => "001000100100111010001",
		474 => "001000111100011110011",
		475 => "001000111100011110011",
		476 => "001000111100011110011",
		477 => "001000100100111010001",
		478 => "001000100100111010001",
		479 => "001000100100111010001",
		480 => "011010100100001010100",
		481 => "011010100100001010100",
		482 => "011010100100001010100",
		483 => "011010100100001010100",
		484 => "011010100100001010100",
		485 => "011010100100001010100",
		486 => "011010100100001010100",
		487 => "011010100100001010100",
		488 => "011010100100001010100",
		489 => "011010100100001010100",
		490 => "011010100100001010100",
		491 => "011010100100001010100",
		492 => "011010100100001010100",
		493 => "011010100100001010100",
		494 => "011010100100001010100",
		495 => "011010100100001010100",
		496 => "011010100100001010100",
		497 => "011010100100001010100",
		498 => "011010100100001010100",
		499 => "011010100100001010100",
		500 => "011010100100001010100",
		501 => "011010100100001010100",
		502 => "011010100100001010100",
		503 => "011010100100001010100",
		504 => "011010100100001010100",
		505 => "011010100100001010100",
		506 => "011010100100001010100",
		507 => "011010100100001010100",
		508 => "011010100100001010100",
		509 => "011010100100001010100",
		510 => "011010100100001010100",
		511 => "011010100100001010100",
		512 => "011010100100001010100",
		513 => "011010100100001010100",
		514 => "011010100100001010100",
		515 => "011010100100001010100",
		516 => "011010100100001010100",
		517 => "011010100100001010100",
		518 => "011010100100001010100",
		519 => "011010100100001010100",
		520 => "011010100100001010100",
		521 => "011010100100001010100",
		522 => "011010100100001010100",
		523 => "011010100100001010100",
		524 => "011010100100001010100",
		525 => "011010100100001010100",
		526 => "011010100100001010100",
		527 => "011010100100001010100",
		528 => "011010100100001010100",
		529 => "011010100100001010100",
		530 => "011010100100001010100",
		531 => "011010100100001010100",
		532 => "011010100100001010100",
		533 => "011010100100001010100",
		534 => "011010100100001010100",
		535 => "011010100100001010100",
		536 => "011010100100001010100",
		537 => "011010100100001010100",
		538 => "011010100100001010100",
		539 => "011010100100001010100",
		540 => "011010100100001010100",
		541 => "011010100100001010100",
		542 => "011010100100001010100",
		543 => "011010100100001010100",
		544 => "011010100100001010100",
		545 => "011010100100001010100",
		546 => "011010100100001010100",
		547 => "011010100100001010100",
		548 => "011010100100001010100",
		549 => "011010100100001010100",
		550 => "011010100100001010100",
		551 => "011010100100001010100",
		552 => "011010100100001010100",
		553 => "011010100100001010100",
		554 => "011010100100001010100",
		555 => "011010100100001010100",
		556 => "011010100100001010100",
		557 => "011010100100001010100",
		558 => "011010100100001010100",
		559 => "011010100100001010100",
		560 => "011010100100001010100",
		561 => "011010100100001010100",
		562 => "011010100100001010100",
		563 => "011010100100001010100",
		564 => "011010100100001010100",
		565 => "011010100100001010100",
		566 => "011010100100001010100",
		567 => "011010100100001010100",
		568 => "011010100100001010100",
		569 => "011010100100001010100",
		570 => "011010100100001010100",
		571 => "011010100100001010100",
		572 => "011010100100001010100",
		573 => "011010100100001010100",
		574 => "011010100100001010100",
		575 => "011010100100001010100",
		576 => "001000111100111010000",
		577 => "001000111100111010000",
		578 => "001000111100111010000",
		579 => "001000111100111010000",
		580 => "001000111100111010000",
		581 => "001000111100111010000",
		582 => "001000111100111010000",
		583 => "001000111100111010000",
		584 => "001000111100111010000",
		585 => "001000111100111010000",
		586 => "001000111100111010000",
		587 => "001000111100111010000",
		588 => "001000111100111010000",
		589 => "001000111100111010000",
		590 => "001000111100111010000",
		591 => "001000111100111010000",
		592 => "001000111100111010000",
		593 => "001000111100111010000",
		594 => "001000111100111010000",
		595 => "001000111100111010000",
		596 => "001000111100111010000",
		597 => "001000111100111010000",
		598 => "001000111100111010000",
		599 => "001000111100111010000",
		600 => "001000111100111010000",
		601 => "001000111100111010000",
		602 => "001000111100111010000",
		603 => "001000111100111010000",
		604 => "001000111100111010000",
		605 => "001000111100111010000",
		606 => "001000111100111010000",
		607 => "001000111100111010000",
		608 => "001000111100111010000",
		609 => "001000111100111010000",
		610 => "001000111100111010000",
		611 => "001000111100111010000",
		612 => "001000111100111010000",
		613 => "001000111100111010000",
		614 => "001000111100111010000",
		615 => "001000111100111010000",
		616 => "001000111100111010000",
		617 => "001000111100111010000",
		618 => "001000111100111010000",
		619 => "001000111100111010000",
		620 => "001000111100111010000",
		621 => "001000111100111010000",
		622 => "001000111100111010000",
		623 => "001000111100111010000",
		624 => "001000111100111010000",
		625 => "001000111100111010000",
		626 => "001000111100111010000",
		627 => "001000111100111010000",
		628 => "001000111100111010000",
		629 => "001000111100111010000",
		630 => "001000111100111010000",
		631 => "001000111100111010000",
		632 => "001000111100111010000",
		633 => "001000111100111010000",
		634 => "001000111100111010000",
		635 => "001000111100111010000",
		636 => "001000111100111010000",
		637 => "001000111100111010000",
		638 => "001000111100111010000",
		639 => "001000111100111010000",
		640 => "001000111100111010000",
		641 => "001000111100111010000",
		642 => "001000111100111010000",
		643 => "001000111100111010000",
		644 => "001000111100111010000",
		645 => "001000111100111010000",
		646 => "001000111100111010000",
		647 => "001000111100111010000",
		648 => "001000111100111010000",
		649 => "001000111100111010000",
		650 => "001000111100111010000",
		651 => "001000111100111010000",
		652 => "001000111100111010000",
		653 => "001000111100111010000",
		654 => "001000111100111010000",
		655 => "001000111100111010000",
		656 => "001000111100111010000",
		657 => "001000111100111010000",
		658 => "001000111100111010000",
		659 => "001000111100111010000",
		660 => "001000111100111010000",
		661 => "001000111100111010000",
		662 => "001000111100111010000",
		663 => "001000111100111010000",
		664 => "001000111100111010000",
		665 => "001000111100111010000",
		666 => "001000111100111010000",
		667 => "001000111100111010000",
		668 => "001000111100111010000",
		669 => "001000111100111010000",
		670 => "001000111100111010000",
		671 => "001000111100111010000",
		672 => "011000101100100010101",
		673 => "011000101100100010101",
		674 => "011000101100100010101",
		675 => "011000101100100010101",
		676 => "011000101100100010101",
		677 => "011000101100100010101",
		678 => "011000101100100010101",
		679 => "011000101100100010101",
		680 => "011000101100100010101",
		681 => "011000101100100010101",
		682 => "011000101100100010101",
		683 => "011000101100100010101",
		684 => "011000101100100010101",
		685 => "011000101100100010101",
		686 => "011000101100100010101",
		687 => "011000101100100010101",
		688 => "011000101100100010101",
		689 => "011000101100100010101",
		690 => "011000101100100010101",
		691 => "011000101100100010101",
		692 => "011000101100100010101",
		693 => "011000101100100010101",
		694 => "011000101100100010101",
		695 => "011000101100100010101",
		696 => "011000101100100010101",
		697 => "011000101100100010101",
		698 => "011000101100100010101",
		699 => "011000101100100010101",
		700 => "011000101100100010101",
		701 => "011000101100100010101",
		702 => "011000101100100010101",
		703 => "011000101100100010101",
		704 => "011000101100100010101",
		705 => "011000101100100010101",
		706 => "011000101100100010101",
		707 => "011000101100100010101",
		708 => "011000101100100010101",
		709 => "011000101100100010101",
		710 => "011000101100100010101",
		711 => "011000101100100010101",
		712 => "011000101100100010101",
		713 => "011000101100100010101",
		714 => "011000101100100010101",
		715 => "011000101100100010101",
		716 => "011000101100100010101",
		717 => "011000101100100010101",
		718 => "011000101100100010101",
		719 => "011000101100100010101",
		720 => "011000101100100010101",
		721 => "011000101100100010101",
		722 => "011000101100100010101",
		723 => "011000101100100010101",
		724 => "011000101100100010101",
		725 => "011000101100100010101",
		726 => "011000101100100010101",
		727 => "011000101100100010101",
		728 => "011000101100100010101",
		729 => "011000101100100010101",
		730 => "011000101100100010101",
		731 => "011000101100100010101",
		732 => "011000101100100010101",
		733 => "011000101100100010101",
		734 => "011000101100100010101",
		735 => "011000101100100010101",
		736 => "011000101100100010101",
		737 => "011000101100100010101",
		738 => "011000101100100010101",
		739 => "011000101100100010101",
		740 => "011000101100100010101",
		741 => "011000101100100010101",
		742 => "011000101100100010101",
		743 => "011000101100100010101",
		744 => "011000101100100010101",
		745 => "011000101100100010101",
		746 => "011000101100100010101",
		747 => "011000101100100010101",
		748 => "011000101100100010101",
		749 => "011000101100100010101",
		750 => "011000101100100010101",
		751 => "011000101100100010101",
		752 => "011000101100100010101",
		753 => "011000101100100010101",
		754 => "011000101100100010101",
		755 => "011000101100100010101",
		756 => "011000101100100010101",
		757 => "011000101100100010101",
		758 => "011000101100100010101",
		759 => "011000101100100010101",
		760 => "011000101100100010101",
		761 => "011000101100100010101",
		762 => "011000101100100010101",
		763 => "011000101100100010101",
		764 => "011000101100100010101",
		765 => "011000101100100010101",
		766 => "011000101100100010101",
		767 => "011000101100100010101",
		768 => "011000101100100110010",
		769 => "011000101100100110010",
		770 => "011000101100100110010",
		771 => "011000101100100110010",
		772 => "011000101100100110010",
		773 => "011000101100100110010",
		774 => "011000101100100110010",
		775 => "011000101100100110010",
		776 => "011000101100100110010",
		777 => "011000101100100110010",
		778 => "011000101100100110010",
		779 => "011000101100100110010",
		780 => "011000101100100110010",
		781 => "011000101100100110010",
		782 => "011000101100100110010",
		783 => "011000101100100110010",
		784 => "011000101100100110010",
		785 => "011000101100100110010",
		786 => "011000101100100110010",
		787 => "011000101100100110010",
		788 => "011000101100100110010",
		789 => "011000101100100110010",
		790 => "011000101100100110010",
		791 => "011000101100100110010",
		792 => "011000101100100110010",
		793 => "011000101100100110010",
		794 => "011000101100100110010",
		795 => "011000101100100110010",
		796 => "011000101100100110010",
		797 => "011000101100100110010",
		798 => "011000101100100110010",
		799 => "011000101100100110010",
		800 => "011000101100100110010",
		801 => "011000101100100110010",
		802 => "011000101100100110010",
		803 => "011000101100100110010",
		804 => "011000101100100110010",
		805 => "011000101100100110010",
		806 => "011000101100100110010",
		807 => "011000101100100110010",
		808 => "011000101100100110010",
		809 => "011000101100100110010",
		810 => "011000101100100110010",
		811 => "011000101100100110010",
		812 => "011000101100100110010",
		813 => "011000101100100110010",
		814 => "011000101100100110010",
		815 => "011000101100100110010",
		816 => "011000101100100110010",
		817 => "011000101100100110010",
		818 => "011000101100100110010",
		819 => "011000101100100110010",
		820 => "011000101100100110010",
		821 => "011000101100100110010",
		822 => "011000101100100110010",
		823 => "011000101100100110010",
		824 => "011000101100100110010",
		825 => "011000101100100110010",
		826 => "011000101100100110010",
		827 => "011000101100100110010",
		828 => "011000101100100110010",
		829 => "011000101100100110010",
		830 => "011000101100100110010",
		831 => "011000101100100110010",
		832 => "011000101100100110010",
		833 => "011000101100100110010",
		834 => "011000101100100110010",
		835 => "011000101100100110010",
		836 => "011000101100100110010",
		837 => "011000101100100110010",
		838 => "011000101100100110010",
		839 => "011000101100100110010",
		840 => "011000101100100110010",
		841 => "011000101100100110010",
		842 => "011000101100100110010",
		843 => "011000101100100110010",
		844 => "011000101100100110010",
		845 => "011000101100100110010",
		846 => "011000101100100110010",
		847 => "011000101100100110010",
		848 => "011000101100100110010",
		849 => "011000101100100110010",
		850 => "011000101100100110010",
		851 => "011000101100100110010",
		852 => "011000101100100110010",
		853 => "011000101100100110010",
		854 => "011000101100100110010",
		855 => "011000101100100110010",
		856 => "011000101100100110010",
		857 => "011000101100100110010",
		858 => "011000101100100110010",
		859 => "011000101100100110010",
		860 => "011000101100100110010",
		861 => "011000101100100110010",
		862 => "011000101100100110010",
		863 => "011000101100100110010");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;