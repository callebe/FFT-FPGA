library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT9 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT9;

architecture Behavioral of ROMFFT9 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 10 
	constant ROM_tb : ROM := (
		0 => "011010011110011010000",
		1 => "011010011110011010000",
		2 => "011010011110011010000",
		3 => "001010111100001110111",
		4 => "001010111100001110111",
		5 => "001010111100001110111",
		6 => "011000000101011110010",
		7 => "011000000101011110010",
		8 => "011000000101011110010",
		9 => "011000111100101010000",
		10 => "011000111100101010000",
		11 => "011000111100101010000",
		12 => "011000001101100010011",
		13 => "011000001101100010011",
		14 => "011000001101100010011",
		15 => "001000011101001010001",
		16 => "001000011101001010001",
		17 => "001000011101001010001",
		18 => "001000111100011110011",
		19 => "001000111100011110011",
		20 => "001000111100011110011",
		21 => "001001011100001010011",
		22 => "001001011100001010011",
		23 => "001001011100001010011",
		24 => "011000101100111010001",
		25 => "011000101100111010001",
		26 => "011000101100111010001",
		27 => "001010011100011110010",
		28 => "001010011100011110010",
		29 => "001010011100011110010",
		30 => "011000111100001010011",
		31 => "011000111100001010011",
		32 => "011000111100001010011",
		33 => "011000001101011010001",
		34 => "011000001101011010001",
		35 => "011000001101011010001",
		36 => "011000011101011010010",
		37 => "011000011101011010010",
		38 => "011000011101011010010",
		39 => "011000001110010010101",
		40 => "011000001110010010101",
		41 => "011000001110010010101",
		42 => "001011011101111010000",
		43 => "001011011101111010000",
		44 => "001011011101111010000",
		45 => "011000000101010011010",
		46 => "011000000101010011010",
		47 => "011000000101010011010",
		48 => "011100100100001010100",
		49 => "011100100100001010100",
		50 => "011100100100001010100",
		51 => "001000000101111010101",
		52 => "001000000101111010101",
		53 => "001000000101111010101",
		54 => "001001011100001010101",
		55 => "001001011100001010101",
		56 => "001001011100001010101",
		57 => "001000111100011110010",
		58 => "001000111100011110010",
		59 => "001000111100011110010",
		60 => "011001100100000010110",
		61 => "011001100100000010110",
		62 => "011001100100000010110",
		63 => "001000011101001010001",
		64 => "001000011101001010001",
		65 => "001000011101001010001",
		66 => "001000100100111010001",
		67 => "001000100100111010001",
		68 => "001000100100111010001",
		69 => "011001100100001010010",
		70 => "011001100100001010010",
		71 => "011001100100001010010",
		72 => "001000110100011010011",
		73 => "001000110100011010011",
		74 => "001000110100011010011",
		75 => "011001000100001010100",
		76 => "011001000100001010100",
		77 => "011001000100001010100",
		78 => "011001100100001110001",
		79 => "011001100100001110001",
		80 => "011001100100001110001",
		81 => "001000000101011110001",
		82 => "001000000101011110001",
		83 => "001000000101011110001",
		84 => "001000011100101010101",
		85 => "001000011100101010101",
		86 => "001000011100101010101",
		87 => "011000001110010010101",
		88 => "011000001110010010101",
		89 => "011000001110010010101",
		90 => "011011100100001110110",
		91 => "011011100100001110110",
		92 => "011011100100001110110",
		93 => "011000000101010011010",
		94 => "011000000101010011010",
		95 => "011000000101010011010",
		96 => "011000000101111010110",
		97 => "011000000101111010110",
		98 => "011000000101111010110",
		99 => "011010100100001010100",
		100 => "011010100100001010100",
		101 => "011010100100001010100",
		102 => "001001011100001010101",
		103 => "001001011100001010101",
		104 => "001001011100001010101",
		105 => "001010111100001110010",
		106 => "001010111100001110010",
		107 => "001010111100001110010",
		108 => "011000101100111010001",
		109 => "011000101100111010001",
		110 => "011000101100111010001",
		111 => "011000000100111010110",
		112 => "011000000100111010110",
		113 => "011000000100111010110",
		114 => "011000000101011010011",
		115 => "011000000101011010011",
		116 => "011000000101011010011",
		117 => "011010111100001011001",
		118 => "011010111100001011001",
		119 => "011010111100001011001",
		120 => "011000000101111010110",
		121 => "011000000101111010110",
		122 => "011000000101111010110",
		123 => "011010100100001010100",
		124 => "011010100100001010100",
		125 => "011010100100001010100",
		126 => "011010100100001010010",
		127 => "011010100100001010010",
		128 => "011010100100001010010",
		129 => "001000000100101010101",
		130 => "001000000100101010101",
		131 => "001000000100101010101",
		132 => "011000101100111010001",
		133 => "011000101100111010001",
		134 => "011000101100111010001",
		135 => "011000000100111010110",
		136 => "011000000100111010110",
		137 => "011000000100111010110",
		138 => "011010100100001110011",
		139 => "011010100100001110011",
		140 => "011010100100001110011",
		141 => "011100100100001110101",
		142 => "011100100100001110101",
		143 => "011100100100001110101",
		144 => "011000000101111010110",
		145 => "011000000101111010110",
		146 => "011000000101111010110",
		147 => "011010100100001010100",
		148 => "011010100100001010100",
		149 => "011010100100001010100",
		150 => "001001011100001010101",
		151 => "001001011100001010101",
		152 => "001001011100001010101",
		153 => "001010111100001110010",
		154 => "001010111100001110010",
		155 => "001010111100001110010",
		156 => "011000101100111010001",
		157 => "011000101100111010001",
		158 => "011000101100111010001",
		159 => "011000000100111010110",
		160 => "011000000100111010110",
		161 => "011000000100111010110",
		162 => "011000000101011010011",
		163 => "011000000101011010011",
		164 => "011000000101011010011",
		165 => "011010111100001011001",
		166 => "011010111100001011001",
		167 => "011010111100001011001",
		168 => "011000000101111010110",
		169 => "011000000101111010110",
		170 => "011000000101111010110",
		171 => "011010100100001010100",
		172 => "011010100100001010100",
		173 => "011010100100001010100",
		174 => "011010100100001010010",
		175 => "011010100100001010010",
		176 => "011010100100001010010",
		177 => "001000000100101010101",
		178 => "001000000100101010101",
		179 => "001000000100101010101",
		180 => "011000101100111010001",
		181 => "011000101100111010001",
		182 => "011000101100111010001",
		183 => "011000000100111010110",
		184 => "011000000100111010110",
		185 => "011000000100111010110",
		186 => "011010100100001110011",
		187 => "011010100100001110011",
		188 => "011010100100001110011",
		189 => "011100100100001110101",
		190 => "011100100100001110101",
		191 => "011100100100001110101",
		192 => "011010100100001010010",
		193 => "011010100100001010010",
		194 => "011010100100001010010",
		195 => "011001111100011110010",
		196 => "011001111100011110010",
		197 => "011001111100011110010",
		198 => "011000000101001010010",
		199 => "011000000101001010010",
		200 => "011000000101001010010",
		201 => "011000000101111010100",
		202 => "011000000101111010100",
		203 => "011000000101111010100",
		204 => "001001011100001010101",
		205 => "001001011100001010101",
		206 => "001001011100001010101",
		207 => "011001000100001110011",
		208 => "011001000100001110011",
		209 => "011001000100001110011",
		210 => "011000000101001010010",
		211 => "011000000101001010010",
		212 => "011000000101001010010",
		213 => "011011100100001110100",
		214 => "011011100100001110100",
		215 => "011011100100001110100",
		216 => "011010100100001010010",
		217 => "011010100100001010010",
		218 => "011010100100001010010",
		219 => "011001111100011110010",
		220 => "011001111100011110010",
		221 => "011001111100011110010",
		222 => "011000000101001010010",
		223 => "011000000101001010010",
		224 => "011000000101001010010",
		225 => "011000000101111010100",
		226 => "011000000101111010100",
		227 => "011000000101111010100",
		228 => "001001011100001010101",
		229 => "001001011100001010101",
		230 => "001001011100001010101",
		231 => "011001000100001110011",
		232 => "011001000100001110011",
		233 => "011001000100001110011",
		234 => "011000000101001010010",
		235 => "011000000101001010010",
		236 => "011000000101001010010",
		237 => "011011100100001110100",
		238 => "011011100100001110100",
		239 => "011011100100001110100",
		240 => "011010100100001010010",
		241 => "011010100100001010010",
		242 => "011010100100001010010",
		243 => "011001111100011110010",
		244 => "011001111100011110010",
		245 => "011001111100011110010",
		246 => "011000000101001010010",
		247 => "011000000101001010010",
		248 => "011000000101001010010",
		249 => "011000000101111010100",
		250 => "011000000101111010100",
		251 => "011000000101111010100",
		252 => "001001011100001010101",
		253 => "001001011100001010101",
		254 => "001001011100001010101",
		255 => "011001000100001110011",
		256 => "011001000100001110011",
		257 => "011001000100001110011",
		258 => "011000000101001010010",
		259 => "011000000101001010010",
		260 => "011000000101001010010",
		261 => "011011100100001110100",
		262 => "011011100100001110100",
		263 => "011011100100001110100",
		264 => "011010100100001010010",
		265 => "011010100100001010010",
		266 => "011010100100001010010",
		267 => "011001111100011110010",
		268 => "011001111100011110010",
		269 => "011001111100011110010",
		270 => "011000000101001010010",
		271 => "011000000101001010010",
		272 => "011000000101001010010",
		273 => "011000000101111010100",
		274 => "011000000101111010100",
		275 => "011000000101111010100",
		276 => "001001011100001010101",
		277 => "001001011100001010101",
		278 => "001001011100001010101",
		279 => "011001000100001110011",
		280 => "011001000100001110011",
		281 => "011001000100001110011",
		282 => "011000000101001010010",
		283 => "011000000101001010010",
		284 => "011000000101001010010",
		285 => "011011100100001110100",
		286 => "011011100100001110100",
		287 => "011011100100001110100",
		288 => "011000000100111010110",
		289 => "011000000100111010110",
		290 => "011000000100111010110",
		291 => "011000000101011010011",
		292 => "011000000101011010011",
		293 => "011000000101011010011",
		294 => "011000001101110010011",
		295 => "011000001101110010011",
		296 => "011000001101110010011",
		297 => "011010100100001110011",
		298 => "011010100100001110011",
		299 => "011010100100001110011",
		300 => "011000000100111010110",
		301 => "011000000100111010110",
		302 => "011000000100111010110",
		303 => "011000000101011010011",
		304 => "011000000101011010011",
		305 => "011000000101011010011",
		306 => "011000001101110010011",
		307 => "011000001101110010011",
		308 => "011000001101110010011",
		309 => "011010100100001110011",
		310 => "011010100100001110011",
		311 => "011010100100001110011",
		312 => "011000000100111010110",
		313 => "011000000100111010110",
		314 => "011000000100111010110",
		315 => "011000000101011010011",
		316 => "011000000101011010011",
		317 => "011000000101011010011",
		318 => "011000001101110010011",
		319 => "011000001101110010011",
		320 => "011000001101110010011",
		321 => "011010100100001110011",
		322 => "011010100100001110011",
		323 => "011010100100001110011",
		324 => "011000000100111010110",
		325 => "011000000100111010110",
		326 => "011000000100111010110",
		327 => "011000000101011010011",
		328 => "011000000101011010011",
		329 => "011000000101011010011",
		330 => "011000001101110010011",
		331 => "011000001101110010011",
		332 => "011000001101110010011",
		333 => "011010100100001110011",
		334 => "011010100100001110011",
		335 => "011010100100001110011",
		336 => "011000000100111010110",
		337 => "011000000100111010110",
		338 => "011000000100111010110",
		339 => "011000000101011010011",
		340 => "011000000101011010011",
		341 => "011000000101011010011",
		342 => "011000001101110010011",
		343 => "011000001101110010011",
		344 => "011000001101110010011",
		345 => "011010100100001110011",
		346 => "011010100100001110011",
		347 => "011010100100001110011",
		348 => "011000000100111010110",
		349 => "011000000100111010110",
		350 => "011000000100111010110",
		351 => "011000000101011010011",
		352 => "011000000101011010011",
		353 => "011000000101011010011",
		354 => "011000001101110010011",
		355 => "011000001101110010011",
		356 => "011000001101110010011",
		357 => "011010100100001110011",
		358 => "011010100100001110011",
		359 => "011010100100001110011",
		360 => "011000000100111010110",
		361 => "011000000100111010110",
		362 => "011000000100111010110",
		363 => "011000000101011010011",
		364 => "011000000101011010011",
		365 => "011000000101011010011",
		366 => "011000001101110010011",
		367 => "011000001101110010011",
		368 => "011000001101110010011",
		369 => "011010100100001110011",
		370 => "011010100100001110011",
		371 => "011010100100001110011",
		372 => "011000000100111010110",
		373 => "011000000100111010110",
		374 => "011000000100111010110",
		375 => "011000000101011010011",
		376 => "011000000101011010011",
		377 => "011000000101011010011",
		378 => "011000001101110010011",
		379 => "011000001101110010011",
		380 => "011000001101110010011",
		381 => "011010100100001110011",
		382 => "011010100100001110011",
		383 => "011010100100001110011",
		384 => "011000101100111010001",
		385 => "011000101100111010001",
		386 => "011000101100111010001",
		387 => "001000000100101110110",
		388 => "001000000100101110110",
		389 => "001000000100101110110",
		390 => "011000101100111010001",
		391 => "011000101100111010001",
		392 => "011000101100111010001",
		393 => "001000000100101110110",
		394 => "001000000100101110110",
		395 => "001000000100101110110",
		396 => "011000101100111010001",
		397 => "011000101100111010001",
		398 => "011000101100111010001",
		399 => "001000000100101110110",
		400 => "001000000100101110110",
		401 => "001000000100101110110",
		402 => "011000101100111010001",
		403 => "011000101100111010001",
		404 => "011000101100111010001",
		405 => "001000000100101110110",
		406 => "001000000100101110110",
		407 => "001000000100101110110",
		408 => "011000101100111010001",
		409 => "011000101100111010001",
		410 => "011000101100111010001",
		411 => "001000000100101110110",
		412 => "001000000100101110110",
		413 => "001000000100101110110",
		414 => "011000101100111010001",
		415 => "011000101100111010001",
		416 => "011000101100111010001",
		417 => "001000000100101110110",
		418 => "001000000100101110110",
		419 => "001000000100101110110",
		420 => "011000101100111010001",
		421 => "011000101100111010001",
		422 => "011000101100111010001",
		423 => "001000000100101110110",
		424 => "001000000100101110110",
		425 => "001000000100101110110",
		426 => "011000101100111010001",
		427 => "011000101100111010001",
		428 => "011000101100111010001",
		429 => "001000000100101110110",
		430 => "001000000100101110110",
		431 => "001000000100101110110",
		432 => "011000101100111010001",
		433 => "011000101100111010001",
		434 => "011000101100111010001",
		435 => "001000000100101110110",
		436 => "001000000100101110110",
		437 => "001000000100101110110",
		438 => "011000101100111010001",
		439 => "011000101100111010001",
		440 => "011000101100111010001",
		441 => "001000000100101110110",
		442 => "001000000100101110110",
		443 => "001000000100101110110",
		444 => "011000101100111010001",
		445 => "011000101100111010001",
		446 => "011000101100111010001",
		447 => "001000000100101110110",
		448 => "001000000100101110110",
		449 => "001000000100101110110",
		450 => "011000101100111010001",
		451 => "011000101100111010001",
		452 => "011000101100111010001",
		453 => "001000000100101110110",
		454 => "001000000100101110110",
		455 => "001000000100101110110",
		456 => "011000101100111010001",
		457 => "011000101100111010001",
		458 => "011000101100111010001",
		459 => "001000000100101110110",
		460 => "001000000100101110110",
		461 => "001000000100101110110",
		462 => "011000101100111010001",
		463 => "011000101100111010001",
		464 => "011000101100111010001",
		465 => "001000000100101110110",
		466 => "001000000100101110110",
		467 => "001000000100101110110",
		468 => "011000101100111010001",
		469 => "011000101100111010001",
		470 => "011000101100111010001",
		471 => "001000000100101110110",
		472 => "001000000100101110110",
		473 => "001000000100101110110",
		474 => "011000101100111010001",
		475 => "011000101100111010001",
		476 => "011000101100111010001",
		477 => "001000000100101110110",
		478 => "001000000100101110110",
		479 => "001000000100101110110",
		480 => "011010100100001110100",
		481 => "011010100100001110100",
		482 => "011010100100001110100",
		483 => "011010100100001110100",
		484 => "011010100100001110100",
		485 => "011010100100001110100",
		486 => "011010100100001110100",
		487 => "011010100100001110100",
		488 => "011010100100001110100",
		489 => "011010100100001110100",
		490 => "011010100100001110100",
		491 => "011010100100001110100",
		492 => "011010100100001110100",
		493 => "011010100100001110100",
		494 => "011010100100001110100",
		495 => "011010100100001110100",
		496 => "011010100100001110100",
		497 => "011010100100001110100",
		498 => "011010100100001110100",
		499 => "011010100100001110100",
		500 => "011010100100001110100",
		501 => "011010100100001110100",
		502 => "011010100100001110100",
		503 => "011010100100001110100",
		504 => "011010100100001110100",
		505 => "011010100100001110100",
		506 => "011010100100001110100",
		507 => "011010100100001110100",
		508 => "011010100100001110100",
		509 => "011010100100001110100",
		510 => "011010100100001110100",
		511 => "011010100100001110100",
		512 => "011010100100001110100",
		513 => "011010100100001110100",
		514 => "011010100100001110100",
		515 => "011010100100001110100",
		516 => "011010100100001110100",
		517 => "011010100100001110100",
		518 => "011010100100001110100",
		519 => "011010100100001110100",
		520 => "011010100100001110100",
		521 => "011010100100001110100",
		522 => "011010100100001110100",
		523 => "011010100100001110100",
		524 => "011010100100001110100",
		525 => "011010100100001110100",
		526 => "011010100100001110100",
		527 => "011010100100001110100",
		528 => "011010100100001110100",
		529 => "011010100100001110100",
		530 => "011010100100001110100",
		531 => "011010100100001110100",
		532 => "011010100100001110100",
		533 => "011010100100001110100",
		534 => "011010100100001110100",
		535 => "011010100100001110100",
		536 => "011010100100001110100",
		537 => "011010100100001110100",
		538 => "011010100100001110100",
		539 => "011010100100001110100",
		540 => "011010100100001110100",
		541 => "011010100100001110100",
		542 => "011010100100001110100",
		543 => "011010100100001110100",
		544 => "011010100100001110100",
		545 => "011010100100001110100",
		546 => "011010100100001110100",
		547 => "011010100100001110100",
		548 => "011010100100001110100",
		549 => "011010100100001110100",
		550 => "011010100100001110100",
		551 => "011010100100001110100",
		552 => "011010100100001110100",
		553 => "011010100100001110100",
		554 => "011010100100001110100",
		555 => "011010100100001110100",
		556 => "011010100100001110100",
		557 => "011010100100001110100",
		558 => "011010100100001110100",
		559 => "011010100100001110100",
		560 => "011010100100001110100",
		561 => "011010100100001110100",
		562 => "011010100100001110100",
		563 => "011010100100001110100",
		564 => "011010100100001110100",
		565 => "011010100100001110100",
		566 => "011010100100001110100",
		567 => "011010100100001110100",
		568 => "011010100100001110100",
		569 => "011010100100001110100",
		570 => "011010100100001110100",
		571 => "011010100100001110100",
		572 => "011010100100001110100",
		573 => "011010100100001110100",
		574 => "011010100100001110100",
		575 => "011010100100001110100",
		576 => "011001111100001010110",
		577 => "011001111100001010110",
		578 => "011001111100001010110",
		579 => "011001111100001010110",
		580 => "011001111100001010110",
		581 => "011001111100001010110",
		582 => "011001111100001010110",
		583 => "011001111100001010110",
		584 => "011001111100001010110",
		585 => "011001111100001010110",
		586 => "011001111100001010110",
		587 => "011001111100001010110",
		588 => "011001111100001010110",
		589 => "011001111100001010110",
		590 => "011001111100001010110",
		591 => "011001111100001010110",
		592 => "011001111100001010110",
		593 => "011001111100001010110",
		594 => "011001111100001010110",
		595 => "011001111100001010110",
		596 => "011001111100001010110",
		597 => "011001111100001010110",
		598 => "011001111100001010110",
		599 => "011001111100001010110",
		600 => "011001111100001010110",
		601 => "011001111100001010110",
		602 => "011001111100001010110",
		603 => "011001111100001010110",
		604 => "011001111100001010110",
		605 => "011001111100001010110",
		606 => "011001111100001010110",
		607 => "011001111100001010110",
		608 => "011001111100001010110",
		609 => "011001111100001010110",
		610 => "011001111100001010110",
		611 => "011001111100001010110",
		612 => "011001111100001010110",
		613 => "011001111100001010110",
		614 => "011001111100001010110",
		615 => "011001111100001010110",
		616 => "011001111100001010110",
		617 => "011001111100001010110",
		618 => "011001111100001010110",
		619 => "011001111100001010110",
		620 => "011001111100001010110",
		621 => "011001111100001010110",
		622 => "011001111100001010110",
		623 => "011001111100001010110",
		624 => "011001111100001010110",
		625 => "011001111100001010110",
		626 => "011001111100001010110",
		627 => "011001111100001010110",
		628 => "011001111100001010110",
		629 => "011001111100001010110",
		630 => "011001111100001010110",
		631 => "011001111100001010110",
		632 => "011001111100001010110",
		633 => "011001111100001010110",
		634 => "011001111100001010110",
		635 => "011001111100001010110",
		636 => "011001111100001010110",
		637 => "011001111100001010110",
		638 => "011001111100001010110",
		639 => "011001111100001010110",
		640 => "011001111100001010110",
		641 => "011001111100001010110",
		642 => "011001111100001010110",
		643 => "011001111100001010110",
		644 => "011001111100001010110",
		645 => "011001111100001010110",
		646 => "011001111100001010110",
		647 => "011001111100001010110",
		648 => "011001111100001010110",
		649 => "011001111100001010110",
		650 => "011001111100001010110",
		651 => "011001111100001010110",
		652 => "011001111100001010110",
		653 => "011001111100001010110",
		654 => "011001111100001010110",
		655 => "011001111100001010110",
		656 => "011001111100001010110",
		657 => "011001111100001010110",
		658 => "011001111100001010110",
		659 => "011001111100001010110",
		660 => "011001111100001010110",
		661 => "011001111100001010110",
		662 => "011001111100001010110",
		663 => "011001111100001010110",
		664 => "011001111100001010110",
		665 => "011001111100001010110",
		666 => "011001111100001010110",
		667 => "011001111100001010110",
		668 => "011001111100001010110",
		669 => "011001111100001010110",
		670 => "011001111100001010110",
		671 => "011001111100001010110",
		672 => "011000101100100010101",
		673 => "011000101100100010101",
		674 => "011000101100100010101",
		675 => "011000101100100010101",
		676 => "011000101100100010101",
		677 => "011000101100100010101",
		678 => "011000101100100010101",
		679 => "011000101100100010101",
		680 => "011000101100100010101",
		681 => "011000101100100010101",
		682 => "011000101100100010101",
		683 => "011000101100100010101",
		684 => "011000101100100010101",
		685 => "011000101100100010101",
		686 => "011000101100100010101",
		687 => "011000101100100010101",
		688 => "011000101100100010101",
		689 => "011000101100100010101",
		690 => "011000101100100010101",
		691 => "011000101100100010101",
		692 => "011000101100100010101",
		693 => "011000101100100010101",
		694 => "011000101100100010101",
		695 => "011000101100100010101",
		696 => "011000101100100010101",
		697 => "011000101100100010101",
		698 => "011000101100100010101",
		699 => "011000101100100010101",
		700 => "011000101100100010101",
		701 => "011000101100100010101",
		702 => "011000101100100010101",
		703 => "011000101100100010101",
		704 => "011000101100100010101",
		705 => "011000101100100010101",
		706 => "011000101100100010101",
		707 => "011000101100100010101",
		708 => "011000101100100010101",
		709 => "011000101100100010101",
		710 => "011000101100100010101",
		711 => "011000101100100010101",
		712 => "011000101100100010101",
		713 => "011000101100100010101",
		714 => "011000101100100010101",
		715 => "011000101100100010101",
		716 => "011000101100100010101",
		717 => "011000101100100010101",
		718 => "011000101100100010101",
		719 => "011000101100100010101",
		720 => "011000101100100010101",
		721 => "011000101100100010101",
		722 => "011000101100100010101",
		723 => "011000101100100010101",
		724 => "011000101100100010101",
		725 => "011000101100100010101",
		726 => "011000101100100010101",
		727 => "011000101100100010101",
		728 => "011000101100100010101",
		729 => "011000101100100010101",
		730 => "011000101100100010101",
		731 => "011000101100100010101",
		732 => "011000101100100010101",
		733 => "011000101100100010101",
		734 => "011000101100100010101",
		735 => "011000101100100010101",
		736 => "011000101100100010101",
		737 => "011000101100100010101",
		738 => "011000101100100010101",
		739 => "011000101100100010101",
		740 => "011000101100100010101",
		741 => "011000101100100010101",
		742 => "011000101100100010101",
		743 => "011000101100100010101",
		744 => "011000101100100010101",
		745 => "011000101100100010101",
		746 => "011000101100100010101",
		747 => "011000101100100010101",
		748 => "011000101100100010101",
		749 => "011000101100100010101",
		750 => "011000101100100010101",
		751 => "011000101100100010101",
		752 => "011000101100100010101",
		753 => "011000101100100010101",
		754 => "011000101100100010101",
		755 => "011000101100100010101",
		756 => "011000101100100010101",
		757 => "011000101100100010101",
		758 => "011000101100100010101",
		759 => "011000101100100010101",
		760 => "011000101100100010101",
		761 => "011000101100100010101",
		762 => "011000101100100010101",
		763 => "011000101100100010101",
		764 => "011000101100100010101",
		765 => "011000101100100010101",
		766 => "011000101100100010101",
		767 => "011000101100100010101",
		768 => "011000101100100110010",
		769 => "011000101100100110010",
		770 => "011000101100100110010",
		771 => "011000101100100110010",
		772 => "011000101100100110010",
		773 => "011000101100100110010",
		774 => "011000101100100110010",
		775 => "011000101100100110010",
		776 => "011000101100100110010",
		777 => "011000101100100110010",
		778 => "011000101100100110010",
		779 => "011000101100100110010",
		780 => "011000101100100110010",
		781 => "011000101100100110010",
		782 => "011000101100100110010",
		783 => "011000101100100110010",
		784 => "011000101100100110010",
		785 => "011000101100100110010",
		786 => "011000101100100110010",
		787 => "011000101100100110010",
		788 => "011000101100100110010",
		789 => "011000101100100110010",
		790 => "011000101100100110010",
		791 => "011000101100100110010",
		792 => "011000101100100110010",
		793 => "011000101100100110010",
		794 => "011000101100100110010",
		795 => "011000101100100110010",
		796 => "011000101100100110010",
		797 => "011000101100100110010",
		798 => "011000101100100110010",
		799 => "011000101100100110010",
		800 => "011000101100100110010",
		801 => "011000101100100110010",
		802 => "011000101100100110010",
		803 => "011000101100100110010",
		804 => "011000101100100110010",
		805 => "011000101100100110010",
		806 => "011000101100100110010",
		807 => "011000101100100110010",
		808 => "011000101100100110010",
		809 => "011000101100100110010",
		810 => "011000101100100110010",
		811 => "011000101100100110010",
		812 => "011000101100100110010",
		813 => "011000101100100110010",
		814 => "011000101100100110010",
		815 => "011000101100100110010",
		816 => "011000101100100110010",
		817 => "011000101100100110010",
		818 => "011000101100100110010",
		819 => "011000101100100110010",
		820 => "011000101100100110010",
		821 => "011000101100100110010",
		822 => "011000101100100110010",
		823 => "011000101100100110010",
		824 => "011000101100100110010",
		825 => "011000101100100110010",
		826 => "011000101100100110010",
		827 => "011000101100100110010",
		828 => "011000101100100110010",
		829 => "011000101100100110010",
		830 => "011000101100100110010",
		831 => "011000101100100110010",
		832 => "011000101100100110010",
		833 => "011000101100100110010",
		834 => "011000101100100110010",
		835 => "011000101100100110010",
		836 => "011000101100100110010",
		837 => "011000101100100110010",
		838 => "011000101100100110010",
		839 => "011000101100100110010",
		840 => "011000101100100110010",
		841 => "011000101100100110010",
		842 => "011000101100100110010",
		843 => "011000101100100110010",
		844 => "011000101100100110010",
		845 => "011000101100100110010",
		846 => "011000101100100110010",
		847 => "011000101100100110010",
		848 => "011000101100100110010",
		849 => "011000101100100110010",
		850 => "011000101100100110010",
		851 => "011000101100100110010",
		852 => "011000101100100110010",
		853 => "011000101100100110010",
		854 => "011000101100100110010",
		855 => "011000101100100110010",
		856 => "011000101100100110010",
		857 => "011000101100100110010",
		858 => "011000101100100110010",
		859 => "011000101100100110010",
		860 => "011000101100100110010",
		861 => "011000101100100110010",
		862 => "011000101100100110010",
		863 => "011000101100100110010");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;