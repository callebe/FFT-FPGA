library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT1024p_2 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT1024p_2;

architecture Behavioral of ROMFFT1024p_2 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 3 
	constant ROM_tb : ROM := (
		0 => "011011000110111010000",
		1 => "011011000110111010000",
		2 => "011011000110111010000",
		3 => "001000011110101010100",
		4 => "001000011110101010100",
		5 => "001000011110101010100",
		6 => "011000000101111010110",
		7 => "011000000101111010110",
		8 => "011000000101111010110",
		9 => "011001111101111010000",
		10 => "011001111101111010000",
		11 => "011001111101111010000",
		12 => "011010100100001110101",
		13 => "011010100100001110101",
		14 => "011010100100001110101",
		15 => "001000010100101011000",
		16 => "001000010100101011000",
		17 => "001000010100101011000",
		18 => "011010100100001010100",
		19 => "011010100100001010100",
		20 => "011010100100001010100",
		21 => "011001001100111010000",
		22 => "011001001100111010000",
		23 => "011001001100111010000",
		24 => "011001011100111010000",
		25 => "011001011100111010000",
		26 => "011001011100111010000",
		27 => "011000001101010010011",
		28 => "011000001101010010011",
		29 => "011000001101010010011",
		30 => "001001011100001010101",
		31 => "001001011100001010101",
		32 => "001001011100001010101",
		33 => "011000111101001010000",
		34 => "011000111101001010000",
		35 => "011000111101001010000",
		36 => "001000111100001110110",
		37 => "001000111100001110110",
		38 => "001000111100001110110",
		39 => "001001111100001010110",
		40 => "001001111100001010110",
		41 => "001001111100001010110",
		42 => "001010111100001110010",
		43 => "001010111100001110010",
		44 => "001010111100001110010",
		45 => "001001011100001010011",
		46 => "001001011100001010011",
		47 => "001001011100001010011",
		48 => "011001100100001110000",
		49 => "011001100100001110000",
		50 => "011001100100001110000",
		51 => "011000000100111110000",
		52 => "011000000100111110000",
		53 => "011000000100111110000",
		54 => "011000101100111010001",
		55 => "011000101100111010001",
		56 => "011000101100111010001",
		57 => "001010011100011110010",
		58 => "001010011100011110010",
		59 => "001010011100011110010",
		60 => "011000010100011010011",
		61 => "011000010100011010011",
		62 => "011000010100011010011",
		63 => "011001100100001110001",
		64 => "011001100100001110001",
		65 => "011001100100001110001",
		66 => "011000000100111010110",
		67 => "011000000100111010110",
		68 => "011000000100111010110",
		69 => "011000000101001010100",
		70 => "011000000101001010100",
		71 => "011000000101001010100",
		72 => "011000001100101010001",
		73 => "011000001100101010001",
		74 => "011000001100101010001",
		75 => "011001100100001110001",
		76 => "011001100100001110001",
		77 => "011001100100001110001",
		78 => "011000000101011010011",
		79 => "011000000101011010011",
		80 => "011000000101011010011",
		81 => "011000000101101010010",
		82 => "011000000101101010010",
		83 => "011000000101101010010",
		84 => "011000000101111010100",
		85 => "011000000101111010100",
		86 => "011000000101111010100",
		87 => "011000000101111010011",
		88 => "011000000101111010011",
		89 => "011000000101111010011",
		90 => "011010111100001011001",
		91 => "011010111100001011001",
		92 => "011010111100001011001",
		93 => "011100001110011110000",
		94 => "011100001110011110000",
		95 => "011100001110011110000",
		96 => "011000000110111110101",
		97 => "011000000110111110101",
		98 => "011000000110111110101",
		99 => "011100000100001010011",
		100 => "011100000100001010011",
		101 => "011100000100001010011",
		102 => "011010100100001010010",
		103 => "011010100100001010010",
		104 => "011010100100001010010",
		105 => "001001011100001010101",
		106 => "001001011100001010101",
		107 => "001001011100001010101",
		108 => "001000111100001110011",
		109 => "001000111100001110011",
		110 => "001000111100001110011",
		111 => "011000000101111011000",
		112 => "011000000101111011000",
		113 => "011000000101111011000",
		114 => "011001111100011110010",
		115 => "011001111100011110010",
		116 => "011001111100011110010",
		117 => "001010011100011110010",
		118 => "001010011100011110010",
		119 => "001010011100011110010",
		120 => "011001100100001110000",
		121 => "011001100100001110000",
		122 => "011001100100001110000",
		123 => "001011011100001110010",
		124 => "001011011100001110010",
		125 => "001011011100001110010",
		126 => "011000000101001010010",
		127 => "011000000101001010010",
		128 => "011000000101001010010",
		129 => "011000001101100010011",
		130 => "011000001101100010011",
		131 => "011000001101100010011",
		132 => "011010100100001110010",
		133 => "011010100100001110010",
		134 => "011010100100001110010",
		135 => "011000000101101010011",
		136 => "011000000101101010011",
		137 => "011000000101101010011",
		138 => "011000000101111010100",
		139 => "011000000101111010100",
		140 => "011000000101111010100",
		141 => "011000011110001010110",
		142 => "011000011110001010110",
		143 => "011000011110001010110",
		144 => "001010111100001011011",
		145 => "001010111100001011011",
		146 => "001010111100001011011",
		147 => "011100000100001111001",
		148 => "011100000100001111001",
		149 => "011100000100001111001",
		150 => "001001011100001010101",
		151 => "001001011100001010101",
		152 => "001001011100001010101",
		153 => "011010100100001010010",
		154 => "011010100100001010010",
		155 => "011010100100001010010",
		156 => "001000111100001110011",
		157 => "001000111100001110011",
		158 => "001000111100001110011",
		159 => "001000111100001010011",
		160 => "001000111100001010011",
		161 => "001000111100001010011",
		162 => "011001000100001110011",
		163 => "011001000100001110011",
		164 => "011001000100001110011",
		165 => "011001000100001010100",
		166 => "011001000100001010100",
		167 => "011001000100001010100",
		168 => "001000011100111010000",
		169 => "001000011100111010000",
		170 => "001000011100111010000",
		171 => "001000000100101010110",
		172 => "001000000100101010110",
		173 => "001000000100101010110",
		174 => "011000000101001010010",
		175 => "011000000101001010010",
		176 => "011000000101001010010",
		177 => "011000001101100010011",
		178 => "011000001101100010011",
		179 => "011000001101100010011",
		180 => "011000000101011010010",
		181 => "011000000101011010010",
		182 => "011000000101011010010",
		183 => "001001100101101010000",
		184 => "001001100101101010000",
		185 => "001001100101101010000",
		186 => "011011100100001110100",
		187 => "011011100100001110100",
		188 => "011011100100001110100",
		189 => "011100000101101010000",
		190 => "011100000101101010000",
		191 => "011100000101101010000",
		192 => "011000000110011110100",
		193 => "011000000110011110100",
		194 => "011000000110011110100",
		195 => "011000001110100010101",
		196 => "011000001110100010101",
		197 => "011000001110100010101",
		198 => "011000000100111010110",
		199 => "011000000100111010110",
		200 => "011000000100111010110",
		201 => "001001111100001010110",
		202 => "001001111100001010110",
		203 => "001001111100001010110",
		204 => "011001011100001010011",
		205 => "011001011100001010011",
		206 => "011001011100001010011",
		207 => "011000111100001010011",
		208 => "011000111100001010011",
		209 => "011000111100001010011",
		210 => "011000000101011010011",
		211 => "011000000101011010011",
		212 => "011000000101011010011",
		213 => "011000010100111010110",
		214 => "011000010100111010110",
		215 => "011000010100111010110",
		216 => "001010011100001011001",
		217 => "001010011100001011001",
		218 => "001010011100001011001",
		219 => "011000001110100010101",
		220 => "011000001110100010101",
		221 => "011000001110100010101",
		222 => "011000001101110010011",
		223 => "011000001101110010011",
		224 => "011000001101110010011",
		225 => "011011000100001010011",
		226 => "011011000100001010011",
		227 => "011011000100001010011",
		228 => "011001100100001110010",
		229 => "011001100100001110010",
		230 => "011001100100001110010",
		231 => "011001100100001110001",
		232 => "011001100100001110001",
		233 => "011001100100001110001",
		234 => "011010100100001110011",
		235 => "011010100100001110011",
		236 => "011010100100001110011",
		237 => "011000000101110011001",
		238 => "011000000101110011001",
		239 => "011000000101110011001",
		240 => "011000000110011110100",
		241 => "011000000110011110100",
		242 => "011000000110011110100",
		243 => "011000001110100010101",
		244 => "011000001110100010101",
		245 => "011000001110100010101",
		246 => "011000000100111010110",
		247 => "011000000100111010110",
		248 => "011000000100111010110",
		249 => "001001111100001010110",
		250 => "001001111100001010110",
		251 => "001001111100001010110",
		252 => "011001011100001010011",
		253 => "011001011100001010011",
		254 => "011001011100001010011",
		255 => "011000111100001010011",
		256 => "011000111100001010011",
		257 => "011000111100001010011",
		258 => "011000000101011010011",
		259 => "011000000101011010011",
		260 => "011000000101011010011",
		261 => "011000010100111010110",
		262 => "011000010100111010110",
		263 => "011000010100111010110",
		264 => "001010011100001011001",
		265 => "001010011100001011001",
		266 => "001010011100001011001",
		267 => "011000001110100010101",
		268 => "011000001110100010101",
		269 => "011000001110100010101",
		270 => "011000001101110010011",
		271 => "011000001101110010011",
		272 => "011000001101110010011",
		273 => "011011000100001010011",
		274 => "011011000100001010011",
		275 => "011011000100001010011",
		276 => "011001100100001110010",
		277 => "011001100100001110010",
		278 => "011001100100001110010",
		279 => "011001100100001110001",
		280 => "011001100100001110001",
		281 => "011001100100001110001",
		282 => "011010100100001110011",
		283 => "011010100100001110011",
		284 => "011010100100001110011",
		285 => "011000000101110011001",
		286 => "011000000101110011001",
		287 => "011000000101110011001",
		288 => "011000000101111110011",
		289 => "011000000101111110011",
		290 => "011000000101111110011",
		291 => "011001011101001010000",
		292 => "011001011101001010000",
		293 => "011001011101001010000",
		294 => "011000101100111010001",
		295 => "011000101100111010001",
		296 => "011000101100111010001",
		297 => "011000000101011010101",
		298 => "011000000101011010101",
		299 => "011000000101011010101",
		300 => "001001111100001010111",
		301 => "001001111100001010111",
		302 => "001001111100001010111",
		303 => "011010000100001010010",
		304 => "011010000100001010010",
		305 => "011010000100001010010",
		306 => "001000000100101110110",
		307 => "001000000100101110110",
		308 => "001000000100101110110",
		309 => "011000000101011010101",
		310 => "011000000101011010101",
		311 => "011000000101011010101",
		312 => "011000000101111110011",
		313 => "011000000101111110011",
		314 => "011000000101111110011",
		315 => "011001011101001010000",
		316 => "011001011101001010000",
		317 => "011001011101001010000",
		318 => "011000101100111010001",
		319 => "011000101100111010001",
		320 => "011000101100111010001",
		321 => "011000000101011010101",
		322 => "011000000101011010101",
		323 => "011000000101011010101",
		324 => "001001111100001010111",
		325 => "001001111100001010111",
		326 => "001001111100001010111",
		327 => "011010000100001010010",
		328 => "011010000100001010010",
		329 => "011010000100001010010",
		330 => "001000000100101110110",
		331 => "001000000100101110110",
		332 => "001000000100101110110",
		333 => "011000000101011010101",
		334 => "011000000101011010101",
		335 => "011000000101011010101",
		336 => "011000000101111110011",
		337 => "011000000101111110011",
		338 => "011000000101111110011",
		339 => "011001011101001010000",
		340 => "011001011101001010000",
		341 => "011001011101001010000",
		342 => "011000101100111010001",
		343 => "011000101100111010001",
		344 => "011000101100111010001",
		345 => "011000000101011010101",
		346 => "011000000101011010101",
		347 => "011000000101011010101",
		348 => "001001111100001010111",
		349 => "001001111100001010111",
		350 => "001001111100001010111",
		351 => "011010000100001010010",
		352 => "011010000100001010010",
		353 => "011010000100001010010",
		354 => "001000000100101110110",
		355 => "001000000100101110110",
		356 => "001000000100101110110",
		357 => "011000000101011010101",
		358 => "011000000101011010101",
		359 => "011000000101011010101",
		360 => "011000000101111110011",
		361 => "011000000101111110011",
		362 => "011000000101111110011",
		363 => "011001011101001010000",
		364 => "011001011101001010000",
		365 => "011001011101001010000",
		366 => "011000101100111010001",
		367 => "011000101100111010001",
		368 => "011000101100111010001",
		369 => "011000000101011010101",
		370 => "011000000101011010101",
		371 => "011000000101011010101",
		372 => "001001111100001010111",
		373 => "001001111100001010111",
		374 => "001001111100001010111",
		375 => "011010000100001010010",
		376 => "011010000100001010010",
		377 => "011010000100001010010",
		378 => "001000000100101110110",
		379 => "001000000100101110110",
		380 => "001000000100101110110",
		381 => "011000000101011010101",
		382 => "011000000101011010101",
		383 => "011000000101011010101",
		384 => "011010100100001110100",
		385 => "011010100100001110100",
		386 => "011010100100001110100",
		387 => "111011010100001010011",
		388 => "111011010100001010011",
		389 => "111011010100001010011",
		390 => "011010100100001110100",
		391 => "011010100100001110100",
		392 => "011010100100001110100",
		393 => "011000001101100010011",
		394 => "011000001101100010011",
		395 => "011000001101100010011",
		396 => "011010100100001110100",
		397 => "011010100100001110100",
		398 => "011010100100001110100",
		399 => "111011010100001010011",
		400 => "111011010100001010011",
		401 => "111011010100001010011",
		402 => "011010100100001110100",
		403 => "011010100100001110100",
		404 => "011010100100001110100",
		405 => "011000001101100010011",
		406 => "011000001101100010011",
		407 => "011000001101100010011",
		408 => "011010100100001110100",
		409 => "011010100100001110100",
		410 => "011010100100001110100",
		411 => "111011010100001010011",
		412 => "111011010100001010011",
		413 => "111011010100001010011",
		414 => "011010100100001110100",
		415 => "011010100100001110100",
		416 => "011010100100001110100",
		417 => "011000001101100010011",
		418 => "011000001101100010011",
		419 => "011000001101100010011",
		420 => "011010100100001110100",
		421 => "011010100100001110100",
		422 => "011010100100001110100",
		423 => "111011010100001010011",
		424 => "111011010100001010011",
		425 => "111011010100001010011",
		426 => "011010100100001110100",
		427 => "011010100100001110100",
		428 => "011010100100001110100",
		429 => "011000001101100010011",
		430 => "011000001101100010011",
		431 => "011000001101100010011",
		432 => "011010100100001110100",
		433 => "011010100100001110100",
		434 => "011010100100001110100",
		435 => "111011010100001010011",
		436 => "111011010100001010011",
		437 => "111011010100001010011",
		438 => "011010100100001110100",
		439 => "011010100100001110100",
		440 => "011010100100001110100",
		441 => "011000001101100010011",
		442 => "011000001101100010011",
		443 => "011000001101100010011",
		444 => "011010100100001110100",
		445 => "011010100100001110100",
		446 => "011010100100001110100",
		447 => "111011010100001010011",
		448 => "111011010100001010011",
		449 => "111011010100001010011",
		450 => "011010100100001110100",
		451 => "011010100100001110100",
		452 => "011010100100001110100",
		453 => "011000001101100010011",
		454 => "011000001101100010011",
		455 => "011000001101100010011",
		456 => "011010100100001110100",
		457 => "011010100100001110100",
		458 => "011010100100001110100",
		459 => "111011010100001010011",
		460 => "111011010100001010011",
		461 => "111011010100001010011",
		462 => "011010100100001110100",
		463 => "011010100100001110100",
		464 => "011010100100001110100",
		465 => "011000001101100010011",
		466 => "011000001101100010011",
		467 => "011000001101100010011",
		468 => "011010100100001110100",
		469 => "011010100100001110100",
		470 => "011010100100001110100",
		471 => "111011010100001010011",
		472 => "111011010100001010011",
		473 => "111011010100001010011",
		474 => "011010100100001110100",
		475 => "011010100100001110100",
		476 => "011010100100001110100",
		477 => "011000001101100010011",
		478 => "011000001101100010011",
		479 => "011000001101100010011",
		480 => "011001111100001010110",
		481 => "011001111100001010110",
		482 => "011001111100001010110",
		483 => "011011000100001110011",
		484 => "011011000100001110011",
		485 => "011011000100001110011",
		486 => "011001111100001010110",
		487 => "011001111100001010110",
		488 => "011001111100001010110",
		489 => "011011000100001110011",
		490 => "011011000100001110011",
		491 => "011011000100001110011",
		492 => "011001111100001010110",
		493 => "011001111100001010110",
		494 => "011001111100001010110",
		495 => "011011000100001110011",
		496 => "011011000100001110011",
		497 => "011011000100001110011",
		498 => "011001111100001010110",
		499 => "011001111100001010110",
		500 => "011001111100001010110",
		501 => "011011000100001110011",
		502 => "011011000100001110011",
		503 => "011011000100001110011",
		504 => "011001111100001010110",
		505 => "011001111100001010110",
		506 => "011001111100001010110",
		507 => "011011000100001110011",
		508 => "011011000100001110011",
		509 => "011011000100001110011",
		510 => "011001111100001010110",
		511 => "011001111100001010110",
		512 => "011001111100001010110",
		513 => "011011000100001110011",
		514 => "011011000100001110011",
		515 => "011011000100001110011",
		516 => "011001111100001010110",
		517 => "011001111100001010110",
		518 => "011001111100001010110",
		519 => "011011000100001110011",
		520 => "011011000100001110011",
		521 => "011011000100001110011",
		522 => "011001111100001010110",
		523 => "011001111100001010110",
		524 => "011001111100001010110",
		525 => "011011000100001110011",
		526 => "011011000100001110011",
		527 => "011011000100001110011",
		528 => "011001111100001010110",
		529 => "011001111100001010110",
		530 => "011001111100001010110",
		531 => "011011000100001110011",
		532 => "011011000100001110011",
		533 => "011011000100001110011",
		534 => "011001111100001010110",
		535 => "011001111100001010110",
		536 => "011001111100001010110",
		537 => "011011000100001110011",
		538 => "011011000100001110011",
		539 => "011011000100001110011",
		540 => "011001111100001010110",
		541 => "011001111100001010110",
		542 => "011001111100001010110",
		543 => "011011000100001110011",
		544 => "011011000100001110011",
		545 => "011011000100001110011",
		546 => "011001111100001010110",
		547 => "011001111100001010110",
		548 => "011001111100001010110",
		549 => "011011000100001110011",
		550 => "011011000100001110011",
		551 => "011011000100001110011",
		552 => "011001111100001010110",
		553 => "011001111100001010110",
		554 => "011001111100001010110",
		555 => "011011000100001110011",
		556 => "011011000100001110011",
		557 => "011011000100001110011",
		558 => "011001111100001010110",
		559 => "011001111100001010110",
		560 => "011001111100001010110",
		561 => "011011000100001110011",
		562 => "011011000100001110011",
		563 => "011011000100001110011",
		564 => "011001111100001010110",
		565 => "011001111100001010110",
		566 => "011001111100001010110",
		567 => "011011000100001110011",
		568 => "011011000100001110011",
		569 => "011011000100001110011",
		570 => "011001111100001010110",
		571 => "011001111100001010110",
		572 => "011001111100001010110",
		573 => "011011000100001110011",
		574 => "011011000100001110011",
		575 => "011011000100001110011",
		576 => "011000101100100010101",
		577 => "011000101100100010101",
		578 => "011000101100100010101",
		579 => "011000101100100010101",
		580 => "011000101100100010101",
		581 => "011000101100100010101",
		582 => "011000101100100010101",
		583 => "011000101100100010101",
		584 => "011000101100100010101",
		585 => "011000101100100010101",
		586 => "011000101100100010101",
		587 => "011000101100100010101",
		588 => "011000101100100010101",
		589 => "011000101100100010101",
		590 => "011000101100100010101",
		591 => "011000101100100010101",
		592 => "011000101100100010101",
		593 => "011000101100100010101",
		594 => "011000101100100010101",
		595 => "011000101100100010101",
		596 => "011000101100100010101",
		597 => "011000101100100010101",
		598 => "011000101100100010101",
		599 => "011000101100100010101",
		600 => "011000101100100010101",
		601 => "011000101100100010101",
		602 => "011000101100100010101",
		603 => "011000101100100010101",
		604 => "011000101100100010101",
		605 => "011000101100100010101",
		606 => "011000101100100010101",
		607 => "011000101100100010101",
		608 => "011000101100100010101",
		609 => "011000101100100010101",
		610 => "011000101100100010101",
		611 => "011000101100100010101",
		612 => "011000101100100010101",
		613 => "011000101100100010101",
		614 => "011000101100100010101",
		615 => "011000101100100010101",
		616 => "011000101100100010101",
		617 => "011000101100100010101",
		618 => "011000101100100010101",
		619 => "011000101100100010101",
		620 => "011000101100100010101",
		621 => "011000101100100010101",
		622 => "011000101100100010101",
		623 => "011000101100100010101",
		624 => "011000101100100010101",
		625 => "011000101100100010101",
		626 => "011000101100100010101",
		627 => "011000101100100010101",
		628 => "011000101100100010101",
		629 => "011000101100100010101",
		630 => "011000101100100010101",
		631 => "011000101100100010101",
		632 => "011000101100100010101",
		633 => "011000101100100010101",
		634 => "011000101100100010101",
		635 => "011000101100100010101",
		636 => "011000101100100010101",
		637 => "011000101100100010101",
		638 => "011000101100100010101",
		639 => "011000101100100010101",
		640 => "011000101100100010101",
		641 => "011000101100100010101",
		642 => "011000101100100010101",
		643 => "011000101100100010101",
		644 => "011000101100100010101",
		645 => "011000101100100010101",
		646 => "011000101100100010101",
		647 => "011000101100100010101",
		648 => "011000101100100010101",
		649 => "011000101100100010101",
		650 => "011000101100100010101",
		651 => "011000101100100010101",
		652 => "011000101100100010101",
		653 => "011000101100100010101",
		654 => "011000101100100010101",
		655 => "011000101100100010101",
		656 => "011000101100100010101",
		657 => "011000101100100010101",
		658 => "011000101100100010101",
		659 => "011000101100100010101",
		660 => "011000101100100010101",
		661 => "011000101100100010101",
		662 => "011000101100100010101",
		663 => "011000101100100010101",
		664 => "011000101100100010101",
		665 => "011000101100100010101",
		666 => "011000101100100010101",
		667 => "011000101100100010101",
		668 => "011000101100100010101",
		669 => "011000101100100010101",
		670 => "011000101100100010101",
		671 => "011000101100100010101",
		672 => "011000101100100110010",
		673 => "011000101100100110010",
		674 => "011000101100100110010",
		675 => "011000101100100110010",
		676 => "011000101100100110010",
		677 => "011000101100100110010",
		678 => "011000101100100110010",
		679 => "011000101100100110010",
		680 => "011000101100100110010",
		681 => "011000101100100110010",
		682 => "011000101100100110010",
		683 => "011000101100100110010",
		684 => "011000101100100110010",
		685 => "011000101100100110010",
		686 => "011000101100100110010",
		687 => "011000101100100110010",
		688 => "011000101100100110010",
		689 => "011000101100100110010",
		690 => "011000101100100110010",
		691 => "011000101100100110010",
		692 => "011000101100100110010",
		693 => "011000101100100110010",
		694 => "011000101100100110010",
		695 => "011000101100100110010",
		696 => "011000101100100110010",
		697 => "011000101100100110010",
		698 => "011000101100100110010",
		699 => "011000101100100110010",
		700 => "011000101100100110010",
		701 => "011000101100100110010",
		702 => "011000101100100110010",
		703 => "011000101100100110010",
		704 => "011000101100100110010",
		705 => "011000101100100110010",
		706 => "011000101100100110010",
		707 => "011000101100100110010",
		708 => "011000101100100110010",
		709 => "011000101100100110010",
		710 => "011000101100100110010",
		711 => "011000101100100110010",
		712 => "011000101100100110010",
		713 => "011000101100100110010",
		714 => "011000101100100110010",
		715 => "011000101100100110010",
		716 => "011000101100100110010",
		717 => "011000101100100110010",
		718 => "011000101100100110010",
		719 => "011000101100100110010",
		720 => "011000101100100110010",
		721 => "011000101100100110010",
		722 => "011000101100100110010",
		723 => "011000101100100110010",
		724 => "011000101100100110010",
		725 => "011000101100100110010",
		726 => "011000101100100110010",
		727 => "011000101100100110010",
		728 => "011000101100100110010",
		729 => "011000101100100110010",
		730 => "011000101100100110010",
		731 => "011000101100100110010",
		732 => "011000101100100110010",
		733 => "011000101100100110010",
		734 => "011000101100100110010",
		735 => "011000101100100110010",
		736 => "011000101100100110010",
		737 => "011000101100100110010",
		738 => "011000101100100110010",
		739 => "011000101100100110010",
		740 => "011000101100100110010",
		741 => "011000101100100110010",
		742 => "011000101100100110010",
		743 => "011000101100100110010",
		744 => "011000101100100110010",
		745 => "011000101100100110010",
		746 => "011000101100100110010",
		747 => "011000101100100110010",
		748 => "011000101100100110010",
		749 => "011000101100100110010",
		750 => "011000101100100110010",
		751 => "011000101100100110010",
		752 => "011000101100100110010",
		753 => "011000101100100110010",
		754 => "011000101100100110010",
		755 => "011000101100100110010",
		756 => "011000101100100110010",
		757 => "011000101100100110010",
		758 => "011000101100100110010",
		759 => "011000101100100110010",
		760 => "011000101100100110010",
		761 => "011000101100100110010",
		762 => "011000101100100110010",
		763 => "011000101100100110010",
		764 => "011000101100100110010",
		765 => "011000101100100110010",
		766 => "011000101100100110010",
		767 => "011000101100100110010",
		768 => "111000010100001010000",
		769 => "111000010100001010000",
		770 => "111000010100001010000",
		771 => "111000010100001010000",
		772 => "111000010100001010000",
		773 => "111000010100001010000",
		774 => "111000010100001010000",
		775 => "111000010100001010000",
		776 => "111000010100001010000",
		777 => "111000010100001010000",
		778 => "111000010100001010000",
		779 => "111000010100001010000",
		780 => "111000010100001010000",
		781 => "111000010100001010000",
		782 => "111000010100001010000",
		783 => "111000010100001010000",
		784 => "111000010100001010000",
		785 => "111000010100001010000",
		786 => "111000010100001010000",
		787 => "111000010100001010000",
		788 => "111000010100001010000",
		789 => "111000010100001010000",
		790 => "111000010100001010000",
		791 => "111000010100001010000",
		792 => "111000010100001010000",
		793 => "111000010100001010000",
		794 => "111000010100001010000",
		795 => "111000010100001010000",
		796 => "111000010100001010000",
		797 => "111000010100001010000",
		798 => "111000010100001010000",
		799 => "111000010100001010000",
		800 => "111000010100001010000",
		801 => "111000010100001010000",
		802 => "111000010100001010000",
		803 => "111000010100001010000",
		804 => "111000010100001010000",
		805 => "111000010100001010000",
		806 => "111000010100001010000",
		807 => "111000010100001010000",
		808 => "111000010100001010000",
		809 => "111000010100001010000",
		810 => "111000010100001010000",
		811 => "111000010100001010000",
		812 => "111000010100001010000",
		813 => "111000010100001010000",
		814 => "111000010100001010000",
		815 => "111000010100001010000",
		816 => "111000010100001010000",
		817 => "111000010100001010000",
		818 => "111000010100001010000",
		819 => "111000010100001010000",
		820 => "111000010100001010000",
		821 => "111000010100001010000",
		822 => "111000010100001010000",
		823 => "111000010100001010000",
		824 => "111000010100001010000",
		825 => "111000010100001010000",
		826 => "111000010100001010000",
		827 => "111000010100001010000",
		828 => "111000010100001010000",
		829 => "111000010100001010000",
		830 => "111000010100001010000",
		831 => "111000010100001010000",
		832 => "111000010100001010000",
		833 => "111000010100001010000",
		834 => "111000010100001010000",
		835 => "111000010100001010000",
		836 => "111000010100001010000",
		837 => "111000010100001010000",
		838 => "111000010100001010000",
		839 => "111000010100001010000",
		840 => "111000010100001010000",
		841 => "111000010100001010000",
		842 => "111000010100001010000",
		843 => "111000010100001010000",
		844 => "111000010100001010000",
		845 => "111000010100001010000",
		846 => "111000010100001010000",
		847 => "111000010100001010000",
		848 => "111000010100001010000",
		849 => "111000010100001010000",
		850 => "111000010100001010000",
		851 => "111000010100001010000",
		852 => "111000010100001010000",
		853 => "111000010100001010000",
		854 => "111000010100001010000",
		855 => "111000010100001010000",
		856 => "111000010100001010000",
		857 => "111000010100001010000",
		858 => "111000010100001010000",
		859 => "111000010100001010000",
		860 => "111000010100001010000",
		861 => "111000010100001010000",
		862 => "111000010100001010000",
		863 => "111000010100001010000");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;