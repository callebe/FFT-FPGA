library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT1024p_1 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT1024p_1;

architecture Behavioral of ROMFFT1024p_1 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 2 
	constant ROM_tb : ROM := (
		0 => "011100100111001110000",
		1 => "011100100111001110000",
		2 => "011100100111001110000",
		3 => "011010011110011010000",
		4 => "011010011110011010000",
		5 => "011010011110011010000",
		6 => "001011011101111010000",
		7 => "001011011101111010000",
		8 => "001011011101111010000",
		9 => "001010111100001110111",
		10 => "001010111100001110111",
		11 => "001010111100001110111",
		12 => "001000010100111010110",
		13 => "001000010100111010110",
		14 => "001000010100111010110",
		15 => "011000000101011110010",
		16 => "011000000101011110010",
		17 => "011000000101011110010",
		18 => "001010011100001010101",
		19 => "001010011100001010101",
		20 => "001010011100001010101",
		21 => "011000111100101010000",
		22 => "011000111100101010000",
		23 => "011000111100101010000",
		24 => "011000111100111010000",
		25 => "011000111100111010000",
		26 => "011000111100111010000",
		27 => "011000001101100010011",
		28 => "011000001101100010011",
		29 => "011000001101100010011",
		30 => "001001011100001010100",
		31 => "001001011100001010100",
		32 => "001001011100001010100",
		33 => "001000011101001010001",
		34 => "001000011101001010001",
		35 => "001000011101001010001",
		36 => "011000001100110010110",
		37 => "011000001100110010110",
		38 => "011000001100110010110",
		39 => "001000111100011110011",
		40 => "001000111100011110011",
		41 => "001000111100011110011",
		42 => "011000101100111110001",
		43 => "011000101100111110001",
		44 => "011000101100111110001",
		45 => "001001011100001010011",
		46 => "001001011100001010011",
		47 => "001001011100001010011",
		48 => "011000000100111010001",
		49 => "011000000100111010001",
		50 => "011000000100111010001",
		51 => "011000101100111010001",
		52 => "011000101100111010001",
		53 => "011000101100111010001",
		54 => "011000101100111010001",
		55 => "011000101100111010001",
		56 => "011000101100111010001",
		57 => "001010011100011110010",
		58 => "001010011100011110010",
		59 => "001010011100011110010",
		60 => "011000000100111010001",
		61 => "011000000100111010001",
		62 => "011000000100111010001",
		63 => "011000111100001010011",
		64 => "011000111100001010011",
		65 => "011000111100001010011",
		66 => "001000111100011110010",
		67 => "001000111100011110010",
		68 => "001000111100011110010",
		69 => "011000001101011010001",
		70 => "011000001101011010001",
		71 => "011000001101011010001",
		72 => "011000000100111010001",
		73 => "011000000100111010001",
		74 => "011000000100111010001",
		75 => "011000011101011010010",
		76 => "011000011101011010010",
		77 => "011000011101011010010",
		78 => "011000000101011010101",
		79 => "011000000101011010101",
		80 => "011000000101011010101",
		81 => "011000001110010010101",
		82 => "011000001110010010101",
		83 => "011000001110010010101",
		84 => "011000000101101010011",
		85 => "011000000101101010011",
		86 => "011000000101101010011",
		87 => "001011011101111010000",
		88 => "001011011101111010000",
		89 => "001011011101111010000",
		90 => "011000000110011010101",
		91 => "011000000110011010101",
		92 => "011000000110011010101",
		93 => "011000000101010011010",
		94 => "011000000101010011010",
		95 => "011000000101010011010",
		96 => "011011000110111010000",
		97 => "011011000110111010000",
		98 => "011011000110111010000",
		99 => "011000000101111010110",
		100 => "011000000101111010110",
		101 => "011000000101111010110",
		102 => "011010100100001110101",
		103 => "011010100100001110101",
		104 => "011010100100001110101",
		105 => "011010100100001010100",
		106 => "011010100100001010100",
		107 => "011010100100001010100",
		108 => "011001011100111010000",
		109 => "011001011100111010000",
		110 => "011001011100111010000",
		111 => "001001011100001010101",
		112 => "001001011100001010101",
		113 => "001001011100001010101",
		114 => "001000111100001110110",
		115 => "001000111100001110110",
		116 => "001000111100001110110",
		117 => "001010111100001110010",
		118 => "001010111100001110010",
		119 => "001010111100001110010",
		120 => "011001100100001110000",
		121 => "011001100100001110000",
		122 => "011001100100001110000",
		123 => "011000101100111010001",
		124 => "011000101100111010001",
		125 => "011000101100111010001",
		126 => "011000010100011010011",
		127 => "011000010100011010011",
		128 => "011000010100011010011",
		129 => "011000000100111010110",
		130 => "011000000100111010110",
		131 => "011000000100111010110",
		132 => "011000001100101010001",
		133 => "011000001100101010001",
		134 => "011000001100101010001",
		135 => "011000000101011010011",
		136 => "011000000101011010011",
		137 => "011000000101011010011",
		138 => "011000000101111010100",
		139 => "011000000101111010100",
		140 => "011000000101111010100",
		141 => "011010111100001011001",
		142 => "011010111100001011001",
		143 => "011010111100001011001",
		144 => "011101100101101110000",
		145 => "011101100101101110000",
		146 => "011101100101101110000",
		147 => "011000000101111010110",
		148 => "011000000101111010110",
		149 => "011000000101111010110",
		150 => "011010100100001110101",
		151 => "011010100100001110101",
		152 => "011010100100001110101",
		153 => "011010100100001010100",
		154 => "011010100100001010100",
		155 => "011010100100001010100",
		156 => "011001011100111010000",
		157 => "011001011100111010000",
		158 => "011001011100111010000",
		159 => "011010100100001010010",
		160 => "011010100100001010010",
		161 => "011010100100001010010",
		162 => "001000000101101010001",
		163 => "001000000101101010001",
		164 => "001000000101101010001",
		165 => "001000000100101010101",
		166 => "001000000100101010101",
		167 => "001000000100101010101",
		168 => "001000011100111010000",
		169 => "001000011100111010000",
		170 => "001000011100111010000",
		171 => "011000101100111010001",
		172 => "011000101100111010001",
		173 => "011000101100111010001",
		174 => "011000010100011010011",
		175 => "011000010100011010011",
		176 => "011000010100011010011",
		177 => "011000000100111010110",
		178 => "011000000100111010110",
		179 => "011000000100111010110",
		180 => "001000000100101110001",
		181 => "001000000100101110001",
		182 => "001000000100101110001",
		183 => "011010100100001110011",
		184 => "011010100100001110011",
		185 => "011010100100001110011",
		186 => "001010011101111010000",
		187 => "001010011101111010000",
		188 => "001010011101111010000",
		189 => "011100100100001110101",
		190 => "011100100100001110101",
		191 => "011100100100001110101",
		192 => "011000000110111110101",
		193 => "011000000110111110101",
		194 => "011000000110111110101",
		195 => "011010100100001010010",
		196 => "011010100100001010010",
		197 => "011010100100001010010",
		198 => "001000111100001110011",
		199 => "001000111100001110011",
		200 => "001000111100001110011",
		201 => "011001111100011110010",
		202 => "011001111100011110010",
		203 => "011001111100011110010",
		204 => "011001100100001110000",
		205 => "011001100100001110000",
		206 => "011001100100001110000",
		207 => "011000000101001010010",
		208 => "011000000101001010010",
		209 => "011000000101001010010",
		210 => "011010100100001110010",
		211 => "011010100100001110010",
		212 => "011010100100001110010",
		213 => "011000000101111010100",
		214 => "011000000101111010100",
		215 => "011000000101111010100",
		216 => "001010111100001011011",
		217 => "001010111100001011011",
		218 => "001010111100001011011",
		219 => "001001011100001010101",
		220 => "001001011100001010101",
		221 => "001001011100001010101",
		222 => "001000111100001110011",
		223 => "001000111100001110011",
		224 => "001000111100001110011",
		225 => "011001000100001110011",
		226 => "011001000100001110011",
		227 => "011001000100001110011",
		228 => "001000011100111010000",
		229 => "001000011100111010000",
		230 => "001000011100111010000",
		231 => "011000000101001010010",
		232 => "011000000101001010010",
		233 => "011000000101001010010",
		234 => "011000000101011010010",
		235 => "011000000101011010010",
		236 => "011000000101011010010",
		237 => "011011100100001110100",
		238 => "011011100100001110100",
		239 => "011011100100001110100",
		240 => "011000000110111110101",
		241 => "011000000110111110101",
		242 => "011000000110111110101",
		243 => "011010100100001010010",
		244 => "011010100100001010010",
		245 => "011010100100001010010",
		246 => "001000111100001110011",
		247 => "001000111100001110011",
		248 => "001000111100001110011",
		249 => "011001111100011110010",
		250 => "011001111100011110010",
		251 => "011001111100011110010",
		252 => "011001100100001110000",
		253 => "011001100100001110000",
		254 => "011001100100001110000",
		255 => "011000000101001010010",
		256 => "011000000101001010010",
		257 => "011000000101001010010",
		258 => "011010100100001110010",
		259 => "011010100100001110010",
		260 => "011010100100001110010",
		261 => "011000000101111010100",
		262 => "011000000101111010100",
		263 => "011000000101111010100",
		264 => "001010111100001011011",
		265 => "001010111100001011011",
		266 => "001010111100001011011",
		267 => "001001011100001010101",
		268 => "001001011100001010101",
		269 => "001001011100001010101",
		270 => "001000111100001110011",
		271 => "001000111100001110011",
		272 => "001000111100001110011",
		273 => "011001000100001110011",
		274 => "011001000100001110011",
		275 => "011001000100001110011",
		276 => "001000011100111010000",
		277 => "001000011100111010000",
		278 => "001000011100111010000",
		279 => "011000000101001010010",
		280 => "011000000101001010010",
		281 => "011000000101001010010",
		282 => "011000000101011010010",
		283 => "011000000101011010010",
		284 => "011000000101011010010",
		285 => "011011100100001110100",
		286 => "011011100100001110100",
		287 => "011011100100001110100",
		288 => "011000000110011110100",
		289 => "011000000110011110100",
		290 => "011000000110011110100",
		291 => "011000000100111010110",
		292 => "011000000100111010110",
		293 => "011000000100111010110",
		294 => "011001011100001010011",
		295 => "011001011100001010011",
		296 => "011001011100001010011",
		297 => "011000000101011010011",
		298 => "011000000101011010011",
		299 => "011000000101011010011",
		300 => "001010011100001011001",
		301 => "001010011100001011001",
		302 => "001010011100001011001",
		303 => "011000001101110010011",
		304 => "011000001101110010011",
		305 => "011000001101110010011",
		306 => "011001100100001110010",
		307 => "011001100100001110010",
		308 => "011001100100001110010",
		309 => "011010100100001110011",
		310 => "011010100100001110011",
		311 => "011010100100001110011",
		312 => "011000000110011110100",
		313 => "011000000110011110100",
		314 => "011000000110011110100",
		315 => "011000000100111010110",
		316 => "011000000100111010110",
		317 => "011000000100111010110",
		318 => "011001011100001010011",
		319 => "011001011100001010011",
		320 => "011001011100001010011",
		321 => "011000000101011010011",
		322 => "011000000101011010011",
		323 => "011000000101011010011",
		324 => "001010011100001011001",
		325 => "001010011100001011001",
		326 => "001010011100001011001",
		327 => "011000001101110010011",
		328 => "011000001101110010011",
		329 => "011000001101110010011",
		330 => "011001100100001110010",
		331 => "011001100100001110010",
		332 => "011001100100001110010",
		333 => "011010100100001110011",
		334 => "011010100100001110011",
		335 => "011010100100001110011",
		336 => "011000000110011110100",
		337 => "011000000110011110100",
		338 => "011000000110011110100",
		339 => "011000000100111010110",
		340 => "011000000100111010110",
		341 => "011000000100111010110",
		342 => "011001011100001010011",
		343 => "011001011100001010011",
		344 => "011001011100001010011",
		345 => "011000000101011010011",
		346 => "011000000101011010011",
		347 => "011000000101011010011",
		348 => "001010011100001011001",
		349 => "001010011100001011001",
		350 => "001010011100001011001",
		351 => "011000001101110010011",
		352 => "011000001101110010011",
		353 => "011000001101110010011",
		354 => "011001100100001110010",
		355 => "011001100100001110010",
		356 => "011001100100001110010",
		357 => "011010100100001110011",
		358 => "011010100100001110011",
		359 => "011010100100001110011",
		360 => "011000000110011110100",
		361 => "011000000110011110100",
		362 => "011000000110011110100",
		363 => "011000000100111010110",
		364 => "011000000100111010110",
		365 => "011000000100111010110",
		366 => "011001011100001010011",
		367 => "011001011100001010011",
		368 => "011001011100001010011",
		369 => "011000000101011010011",
		370 => "011000000101011010011",
		371 => "011000000101011010011",
		372 => "001010011100001011001",
		373 => "001010011100001011001",
		374 => "001010011100001011001",
		375 => "011000001101110010011",
		376 => "011000001101110010011",
		377 => "011000001101110010011",
		378 => "011001100100001110010",
		379 => "011001100100001110010",
		380 => "011001100100001110010",
		381 => "011010100100001110011",
		382 => "011010100100001110011",
		383 => "011010100100001110011",
		384 => "011000000101111110011",
		385 => "011000000101111110011",
		386 => "011000000101111110011",
		387 => "011000101100111010001",
		388 => "011000101100111010001",
		389 => "011000101100111010001",
		390 => "001001111100001010111",
		391 => "001001111100001010111",
		392 => "001001111100001010111",
		393 => "001000000100101110110",
		394 => "001000000100101110110",
		395 => "001000000100101110110",
		396 => "011000000101111110011",
		397 => "011000000101111110011",
		398 => "011000000101111110011",
		399 => "011000101100111010001",
		400 => "011000101100111010001",
		401 => "011000101100111010001",
		402 => "001001111100001010111",
		403 => "001001111100001010111",
		404 => "001001111100001010111",
		405 => "001000000100101110110",
		406 => "001000000100101110110",
		407 => "001000000100101110110",
		408 => "011000000101111110011",
		409 => "011000000101111110011",
		410 => "011000000101111110011",
		411 => "011000101100111010001",
		412 => "011000101100111010001",
		413 => "011000101100111010001",
		414 => "001001111100001010111",
		415 => "001001111100001010111",
		416 => "001001111100001010111",
		417 => "001000000100101110110",
		418 => "001000000100101110110",
		419 => "001000000100101110110",
		420 => "011000000101111110011",
		421 => "011000000101111110011",
		422 => "011000000101111110011",
		423 => "011000101100111010001",
		424 => "011000101100111010001",
		425 => "011000101100111010001",
		426 => "001001111100001010111",
		427 => "001001111100001010111",
		428 => "001001111100001010111",
		429 => "001000000100101110110",
		430 => "001000000100101110110",
		431 => "001000000100101110110",
		432 => "011000000101111110011",
		433 => "011000000101111110011",
		434 => "011000000101111110011",
		435 => "011000101100111010001",
		436 => "011000101100111010001",
		437 => "011000101100111010001",
		438 => "001001111100001010111",
		439 => "001001111100001010111",
		440 => "001001111100001010111",
		441 => "001000000100101110110",
		442 => "001000000100101110110",
		443 => "001000000100101110110",
		444 => "011000000101111110011",
		445 => "011000000101111110011",
		446 => "011000000101111110011",
		447 => "011000101100111010001",
		448 => "011000101100111010001",
		449 => "011000101100111010001",
		450 => "001001111100001010111",
		451 => "001001111100001010111",
		452 => "001001111100001010111",
		453 => "001000000100101110110",
		454 => "001000000100101110110",
		455 => "001000000100101110110",
		456 => "011000000101111110011",
		457 => "011000000101111110011",
		458 => "011000000101111110011",
		459 => "011000101100111010001",
		460 => "011000101100111010001",
		461 => "011000101100111010001",
		462 => "001001111100001010111",
		463 => "001001111100001010111",
		464 => "001001111100001010111",
		465 => "001000000100101110110",
		466 => "001000000100101110110",
		467 => "001000000100101110110",
		468 => "011000000101111110011",
		469 => "011000000101111110011",
		470 => "011000000101111110011",
		471 => "011000101100111010001",
		472 => "011000101100111010001",
		473 => "011000101100111010001",
		474 => "001001111100001010111",
		475 => "001001111100001010111",
		476 => "001001111100001010111",
		477 => "001000000100101110110",
		478 => "001000000100101110110",
		479 => "001000000100101110110",
		480 => "011010100100001110100",
		481 => "011010100100001110100",
		482 => "011010100100001110100",
		483 => "011010100100001110100",
		484 => "011010100100001110100",
		485 => "011010100100001110100",
		486 => "011010100100001110100",
		487 => "011010100100001110100",
		488 => "011010100100001110100",
		489 => "011010100100001110100",
		490 => "011010100100001110100",
		491 => "011010100100001110100",
		492 => "011010100100001110100",
		493 => "011010100100001110100",
		494 => "011010100100001110100",
		495 => "011010100100001110100",
		496 => "011010100100001110100",
		497 => "011010100100001110100",
		498 => "011010100100001110100",
		499 => "011010100100001110100",
		500 => "011010100100001110100",
		501 => "011010100100001110100",
		502 => "011010100100001110100",
		503 => "011010100100001110100",
		504 => "011010100100001110100",
		505 => "011010100100001110100",
		506 => "011010100100001110100",
		507 => "011010100100001110100",
		508 => "011010100100001110100",
		509 => "011010100100001110100",
		510 => "011010100100001110100",
		511 => "011010100100001110100",
		512 => "011010100100001110100",
		513 => "011010100100001110100",
		514 => "011010100100001110100",
		515 => "011010100100001110100",
		516 => "011010100100001110100",
		517 => "011010100100001110100",
		518 => "011010100100001110100",
		519 => "011010100100001110100",
		520 => "011010100100001110100",
		521 => "011010100100001110100",
		522 => "011010100100001110100",
		523 => "011010100100001110100",
		524 => "011010100100001110100",
		525 => "011010100100001110100",
		526 => "011010100100001110100",
		527 => "011010100100001110100",
		528 => "011010100100001110100",
		529 => "011010100100001110100",
		530 => "011010100100001110100",
		531 => "011010100100001110100",
		532 => "011010100100001110100",
		533 => "011010100100001110100",
		534 => "011010100100001110100",
		535 => "011010100100001110100",
		536 => "011010100100001110100",
		537 => "011010100100001110100",
		538 => "011010100100001110100",
		539 => "011010100100001110100",
		540 => "011010100100001110100",
		541 => "011010100100001110100",
		542 => "011010100100001110100",
		543 => "011010100100001110100",
		544 => "011010100100001110100",
		545 => "011010100100001110100",
		546 => "011010100100001110100",
		547 => "011010100100001110100",
		548 => "011010100100001110100",
		549 => "011010100100001110100",
		550 => "011010100100001110100",
		551 => "011010100100001110100",
		552 => "011010100100001110100",
		553 => "011010100100001110100",
		554 => "011010100100001110100",
		555 => "011010100100001110100",
		556 => "011010100100001110100",
		557 => "011010100100001110100",
		558 => "011010100100001110100",
		559 => "011010100100001110100",
		560 => "011010100100001110100",
		561 => "011010100100001110100",
		562 => "011010100100001110100",
		563 => "011010100100001110100",
		564 => "011010100100001110100",
		565 => "011010100100001110100",
		566 => "011010100100001110100",
		567 => "011010100100001110100",
		568 => "011010100100001110100",
		569 => "011010100100001110100",
		570 => "011010100100001110100",
		571 => "011010100100001110100",
		572 => "011010100100001110100",
		573 => "011010100100001110100",
		574 => "011010100100001110100",
		575 => "011010100100001110100",
		576 => "011001111100001010110",
		577 => "011001111100001010110",
		578 => "011001111100001010110",
		579 => "011001111100001010110",
		580 => "011001111100001010110",
		581 => "011001111100001010110",
		582 => "011001111100001010110",
		583 => "011001111100001010110",
		584 => "011001111100001010110",
		585 => "011001111100001010110",
		586 => "011001111100001010110",
		587 => "011001111100001010110",
		588 => "011001111100001010110",
		589 => "011001111100001010110",
		590 => "011001111100001010110",
		591 => "011001111100001010110",
		592 => "011001111100001010110",
		593 => "011001111100001010110",
		594 => "011001111100001010110",
		595 => "011001111100001010110",
		596 => "011001111100001010110",
		597 => "011001111100001010110",
		598 => "011001111100001010110",
		599 => "011001111100001010110",
		600 => "011001111100001010110",
		601 => "011001111100001010110",
		602 => "011001111100001010110",
		603 => "011001111100001010110",
		604 => "011001111100001010110",
		605 => "011001111100001010110",
		606 => "011001111100001010110",
		607 => "011001111100001010110",
		608 => "011001111100001010110",
		609 => "011001111100001010110",
		610 => "011001111100001010110",
		611 => "011001111100001010110",
		612 => "011001111100001010110",
		613 => "011001111100001010110",
		614 => "011001111100001010110",
		615 => "011001111100001010110",
		616 => "011001111100001010110",
		617 => "011001111100001010110",
		618 => "011001111100001010110",
		619 => "011001111100001010110",
		620 => "011001111100001010110",
		621 => "011001111100001010110",
		622 => "011001111100001010110",
		623 => "011001111100001010110",
		624 => "011001111100001010110",
		625 => "011001111100001010110",
		626 => "011001111100001010110",
		627 => "011001111100001010110",
		628 => "011001111100001010110",
		629 => "011001111100001010110",
		630 => "011001111100001010110",
		631 => "011001111100001010110",
		632 => "011001111100001010110",
		633 => "011001111100001010110",
		634 => "011001111100001010110",
		635 => "011001111100001010110",
		636 => "011001111100001010110",
		637 => "011001111100001010110",
		638 => "011001111100001010110",
		639 => "011001111100001010110",
		640 => "011001111100001010110",
		641 => "011001111100001010110",
		642 => "011001111100001010110",
		643 => "011001111100001010110",
		644 => "011001111100001010110",
		645 => "011001111100001010110",
		646 => "011001111100001010110",
		647 => "011001111100001010110",
		648 => "011001111100001010110",
		649 => "011001111100001010110",
		650 => "011001111100001010110",
		651 => "011001111100001010110",
		652 => "011001111100001010110",
		653 => "011001111100001010110",
		654 => "011001111100001010110",
		655 => "011001111100001010110",
		656 => "011001111100001010110",
		657 => "011001111100001010110",
		658 => "011001111100001010110",
		659 => "011001111100001010110",
		660 => "011001111100001010110",
		661 => "011001111100001010110",
		662 => "011001111100001010110",
		663 => "011001111100001010110",
		664 => "011001111100001010110",
		665 => "011001111100001010110",
		666 => "011001111100001010110",
		667 => "011001111100001010110",
		668 => "011001111100001010110",
		669 => "011001111100001010110",
		670 => "011001111100001010110",
		671 => "011001111100001010110",
		672 => "011000101100100010101",
		673 => "011000101100100010101",
		674 => "011000101100100010101",
		675 => "011000101100100010101",
		676 => "011000101100100010101",
		677 => "011000101100100010101",
		678 => "011000101100100010101",
		679 => "011000101100100010101",
		680 => "011000101100100010101",
		681 => "011000101100100010101",
		682 => "011000101100100010101",
		683 => "011000101100100010101",
		684 => "011000101100100010101",
		685 => "011000101100100010101",
		686 => "011000101100100010101",
		687 => "011000101100100010101",
		688 => "011000101100100010101",
		689 => "011000101100100010101",
		690 => "011000101100100010101",
		691 => "011000101100100010101",
		692 => "011000101100100010101",
		693 => "011000101100100010101",
		694 => "011000101100100010101",
		695 => "011000101100100010101",
		696 => "011000101100100010101",
		697 => "011000101100100010101",
		698 => "011000101100100010101",
		699 => "011000101100100010101",
		700 => "011000101100100010101",
		701 => "011000101100100010101",
		702 => "011000101100100010101",
		703 => "011000101100100010101",
		704 => "011000101100100010101",
		705 => "011000101100100010101",
		706 => "011000101100100010101",
		707 => "011000101100100010101",
		708 => "011000101100100010101",
		709 => "011000101100100010101",
		710 => "011000101100100010101",
		711 => "011000101100100010101",
		712 => "011000101100100010101",
		713 => "011000101100100010101",
		714 => "011000101100100010101",
		715 => "011000101100100010101",
		716 => "011000101100100010101",
		717 => "011000101100100010101",
		718 => "011000101100100010101",
		719 => "011000101100100010101",
		720 => "011000101100100010101",
		721 => "011000101100100010101",
		722 => "011000101100100010101",
		723 => "011000101100100010101",
		724 => "011000101100100010101",
		725 => "011000101100100010101",
		726 => "011000101100100010101",
		727 => "011000101100100010101",
		728 => "011000101100100010101",
		729 => "011000101100100010101",
		730 => "011000101100100010101",
		731 => "011000101100100010101",
		732 => "011000101100100010101",
		733 => "011000101100100010101",
		734 => "011000101100100010101",
		735 => "011000101100100010101",
		736 => "011000101100100010101",
		737 => "011000101100100010101",
		738 => "011000101100100010101",
		739 => "011000101100100010101",
		740 => "011000101100100010101",
		741 => "011000101100100010101",
		742 => "011000101100100010101",
		743 => "011000101100100010101",
		744 => "011000101100100010101",
		745 => "011000101100100010101",
		746 => "011000101100100010101",
		747 => "011000101100100010101",
		748 => "011000101100100010101",
		749 => "011000101100100010101",
		750 => "011000101100100010101",
		751 => "011000101100100010101",
		752 => "011000101100100010101",
		753 => "011000101100100010101",
		754 => "011000101100100010101",
		755 => "011000101100100010101",
		756 => "011000101100100010101",
		757 => "011000101100100010101",
		758 => "011000101100100010101",
		759 => "011000101100100010101",
		760 => "011000101100100010101",
		761 => "011000101100100010101",
		762 => "011000101100100010101",
		763 => "011000101100100010101",
		764 => "011000101100100010101",
		765 => "011000101100100010101",
		766 => "011000101100100010101",
		767 => "011000101100100010101",
		768 => "011000101100100110010",
		769 => "011000101100100110010",
		770 => "011000101100100110010",
		771 => "011000101100100110010",
		772 => "011000101100100110010",
		773 => "011000101100100110010",
		774 => "011000101100100110010",
		775 => "011000101100100110010",
		776 => "011000101100100110010",
		777 => "011000101100100110010",
		778 => "011000101100100110010",
		779 => "011000101100100110010",
		780 => "011000101100100110010",
		781 => "011000101100100110010",
		782 => "011000101100100110010",
		783 => "011000101100100110010",
		784 => "011000101100100110010",
		785 => "011000101100100110010",
		786 => "011000101100100110010",
		787 => "011000101100100110010",
		788 => "011000101100100110010",
		789 => "011000101100100110010",
		790 => "011000101100100110010",
		791 => "011000101100100110010",
		792 => "011000101100100110010",
		793 => "011000101100100110010",
		794 => "011000101100100110010",
		795 => "011000101100100110010",
		796 => "011000101100100110010",
		797 => "011000101100100110010",
		798 => "011000101100100110010",
		799 => "011000101100100110010",
		800 => "011000101100100110010",
		801 => "011000101100100110010",
		802 => "011000101100100110010",
		803 => "011000101100100110010",
		804 => "011000101100100110010",
		805 => "011000101100100110010",
		806 => "011000101100100110010",
		807 => "011000101100100110010",
		808 => "011000101100100110010",
		809 => "011000101100100110010",
		810 => "011000101100100110010",
		811 => "011000101100100110010",
		812 => "011000101100100110010",
		813 => "011000101100100110010",
		814 => "011000101100100110010",
		815 => "011000101100100110010",
		816 => "011000101100100110010",
		817 => "011000101100100110010",
		818 => "011000101100100110010",
		819 => "011000101100100110010",
		820 => "011000101100100110010",
		821 => "011000101100100110010",
		822 => "011000101100100110010",
		823 => "011000101100100110010",
		824 => "011000101100100110010",
		825 => "011000101100100110010",
		826 => "011000101100100110010",
		827 => "011000101100100110010",
		828 => "011000101100100110010",
		829 => "011000101100100110010",
		830 => "011000101100100110010",
		831 => "011000101100100110010",
		832 => "011000101100100110010",
		833 => "011000101100100110010",
		834 => "011000101100100110010",
		835 => "011000101100100110010",
		836 => "011000101100100110010",
		837 => "011000101100100110010",
		838 => "011000101100100110010",
		839 => "011000101100100110010",
		840 => "011000101100100110010",
		841 => "011000101100100110010",
		842 => "011000101100100110010",
		843 => "011000101100100110010",
		844 => "011000101100100110010",
		845 => "011000101100100110010",
		846 => "011000101100100110010",
		847 => "011000101100100110010",
		848 => "011000101100100110010",
		849 => "011000101100100110010",
		850 => "011000101100100110010",
		851 => "011000101100100110010",
		852 => "011000101100100110010",
		853 => "011000101100100110010",
		854 => "011000101100100110010",
		855 => "011000101100100110010",
		856 => "011000101100100110010",
		857 => "011000101100100110010",
		858 => "011000101100100110010",
		859 => "011000101100100110010",
		860 => "011000101100100110010",
		861 => "011000101100100110010",
		862 => "011000101100100110010",
		863 => "011000101100100110010");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;