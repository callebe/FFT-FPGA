library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT1024p_0 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT1024p_0;

architecture Behavioral of ROMFFT1024p_0 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 1 
	constant ROM_tb : ROM := (
		0 => "111000010100001010000",
		1 => "111000010100001010000",
		2 => "111000010100001010000",
		3 => "011000000110011110100",
		4 => "011000000110011110100",
		5 => "011000000110011110100",
		6 => "011000000101111110011",
		7 => "011000000101111110011",
		8 => "011000000101111110011",
		9 => "011000000101110011001",
		10 => "011000000101110011001",
		11 => "011000000101110011001",
		12 => "011010100100001110100",
		13 => "011010100100001110100",
		14 => "011010100100001110100",
		15 => "011000001110100010101",
		16 => "011000001110100010101",
		17 => "011000001110100010101",
		18 => "001010111100001010101",
		19 => "001010111100001010101",
		20 => "001010111100001010101",
		21 => "001001111100001010101",
		22 => "001001111100001010101",
		23 => "001001111100001010101",
		24 => "011001111100001010110",
		25 => "011001111100001010110",
		26 => "011001111100001010110",
		27 => "011000000100111010110",
		28 => "011000000100111010110",
		29 => "011000000100111010110",
		30 => "011001011101001010000",
		31 => "011001011101001010000",
		32 => "011001011101001010000",
		33 => "001011011100001010111",
		34 => "001011011100001010111",
		35 => "001011011100001010111",
		36 => "011000001101100010011",
		37 => "011000001101100010011",
		38 => "011000001101100010011",
		39 => "001001111100001010110",
		40 => "001001111100001010110",
		41 => "001001111100001010110",
		42 => "001000111100011110011",
		43 => "001000111100011110011",
		44 => "001000111100011110011",
		45 => "011001011100111010000",
		46 => "011001011100111010000",
		47 => "011001011100111010000",
		48 => "011000101100100010101",
		49 => "011000101100100010101",
		50 => "011000101100100010101",
		51 => "011001011100001010011",
		52 => "011001011100001010011",
		53 => "011001011100001010011",
		54 => "011000101100111010001",
		55 => "011000101100111010001",
		56 => "011000101100111010001",
		57 => "011000000101101010011",
		58 => "011000000101101010011",
		59 => "011000000101101010011",
		60 => "111011010100001010011",
		61 => "111011010100001010011",
		62 => "111011010100001010011",
		63 => "011000111100001010011",
		64 => "011000111100001010011",
		65 => "011000111100001010011",
		66 => "011001011100001010100",
		67 => "011001011100001010100",
		68 => "011001011100001010100",
		69 => "011000001101110010011",
		70 => "011000001101110010011",
		71 => "011000001101110010011",
		72 => "011001100100001110001",
		73 => "011001100100001110001",
		74 => "011001100100001110001",
		75 => "011000000101011010011",
		76 => "011000000101011010011",
		77 => "011000000101011010011",
		78 => "011000000101011010101",
		79 => "011000000101011010101",
		80 => "011000000101011010101",
		81 => "011000001110100010101",
		82 => "011000001110100010101",
		83 => "011000001110100010101",
		84 => "011010100100001010100",
		85 => "011010100100001010100",
		86 => "011010100100001010100",
		87 => "011000010100111010110",
		88 => "011000010100111010110",
		89 => "011000010100111010110",
		90 => "011011100100001110011",
		91 => "011011100100001110011",
		92 => "011011100100001110011",
		93 => "011000000110011010100",
		94 => "011000000110011010100",
		95 => "011000000110011010100",
		96 => "011000101100100110010",
		97 => "011000101100100110010",
		98 => "011000101100100110010",
		99 => "001010011100001011001",
		100 => "001010011100001011001",
		101 => "001010011100001011001",
		102 => "001001111100001010111",
		103 => "001001111100001010111",
		104 => "001001111100001010111",
		105 => "011000000101110011001",
		106 => "011000000101110011001",
		107 => "011000000101110011001",
		108 => "011010100100001110100",
		109 => "011010100100001110100",
		110 => "011010100100001110100",
		111 => "011000001110100010101",
		112 => "011000001110100010101",
		113 => "011000001110100010101",
		114 => "011010100100001010101",
		115 => "011010100100001010101",
		116 => "011010100100001010101",
		117 => "001000011101011010010",
		118 => "001000011101011010010",
		119 => "001000011101011010010",
		120 => "011011000100001110011",
		121 => "011011000100001110011",
		122 => "011011000100001110011",
		123 => "011000001101110010011",
		124 => "011000001101110010011",
		125 => "011000001101110010011",
		126 => "011010000100001010010",
		127 => "011010000100001010010",
		128 => "011010000100001010010",
		129 => "011000111100111010000",
		130 => "011000111100111010000",
		131 => "011000111100111010000",
		132 => "011000001101100010011",
		133 => "011000001101100010011",
		134 => "011000001101100010011",
		135 => "011011000100001010011",
		136 => "011011000100001010011",
		137 => "011011000100001010011",
		138 => "001000100100111010001",
		139 => "001000100100111010001",
		140 => "001000100100111010001",
		141 => "011001100100001010010",
		142 => "011001100100001010010",
		143 => "011001100100001010010",
		144 => "011000101100100010101",
		145 => "011000101100100010101",
		146 => "011000101100100010101",
		147 => "011001100100001110010",
		148 => "011001100100001110010",
		149 => "011001100100001110010",
		150 => "001000000100101110110",
		151 => "001000000100101110110",
		152 => "001000000100101110110",
		153 => "011000000101101010011",
		154 => "011000000101101010011",
		155 => "011000000101101010011",
		156 => "011000001101100010011",
		157 => "011000001101100010011",
		158 => "011000001101100010011",
		159 => "011001100100001110001",
		160 => "011001100100001110001",
		161 => "011001100100001110001",
		162 => "011010000100001110010",
		163 => "011010000100001110010",
		164 => "011010000100001110010",
		165 => "011000001101110010011",
		166 => "011000001101110010011",
		167 => "011000001101110010011",
		168 => "001000111100111010000",
		169 => "001000111100111010000",
		170 => "001000111100111010000",
		171 => "011010100100001110011",
		172 => "011010100100001110011",
		173 => "011010100100001110011",
		174 => "011000000101011010101",
		175 => "011000000101011010101",
		176 => "011000000101011010101",
		177 => "011000001110100010101",
		178 => "011000001110100010101",
		179 => "011000001110100010101",
		180 => "011010100100001010100",
		181 => "011010100100001010100",
		182 => "011010100100001010100",
		183 => "011000000101110011001",
		184 => "011000000101110011001",
		185 => "011000000101110011001",
		186 => "011000000101111010011",
		187 => "011000000101111010011",
		188 => "011000000101111010011",
		189 => "001010011110011010000",
		190 => "001010011110011010000",
		191 => "001010011110011010000",
