library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT11 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT11;

architecture Behavioral of ROMFFT11 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 12 
	constant ROM_tb : ROM := (
		0 => "011100011110011010000",
		1 => "011100011110011010000",
		2 => "011100011110011010000",
		3 => "011001111100101010000",
		4 => "011001111100101010000",
		5 => "011001111100101010000",
		6 => "011000000101101110010",
		7 => "011000000101101110010",
		8 => "011000000101101110010",
		9 => "011000000100111010011",
		10 => "011000000100111010011",
		11 => "011000000100111010011",
		12 => "011000000100111010110",
		13 => "011000000100111010110",
		14 => "011000000100111010110",
		15 => "001000111100001010011",
		16 => "001000111100001010011",
		17 => "001000111100001010011",
		18 => "011000000100111010000",
		19 => "011000000100111010000",
		20 => "011000000100111010000",
		21 => "001001011100001010011",
		22 => "001001011100001010011",
		23 => "001001011100001010011",
		24 => "011000011100111010000",
		25 => "011000011100111010000",
		26 => "011000011100111010000",
		27 => "001001111100011110010",
		28 => "001001111100011110010",
		29 => "001001111100011110010",
		30 => "011000000100111010001",
		31 => "011000000100111010001",
		32 => "011000000100111010001",
		33 => "011010000100001110001",
		34 => "011010000100001110001",
		35 => "011010000100001110001",
		36 => "011000000101011010100",
		37 => "011000000101011010100",
		38 => "011000000101011010100",
		39 => "011011011101011010000",
		40 => "011011011101011010000",
		41 => "011011011101011010000",
		42 => "011000010101001011000",
		43 => "011000010101001011000",
		44 => "011000010101001011000",
		45 => "011101100100001011011",
		46 => "011101100100001011011",
		47 => "011101100100001011011",
		48 => "011100100100001011000",
		49 => "011100100100001011000",
		50 => "011100100100001011000",
		51 => "011000001100100110100",
		52 => "011000001100100110100",
		53 => "011000001100100110100",
		54 => "001001011100001010110",
		55 => "001001011100001010110",
		56 => "001001011100001010110",
		57 => "011001100100001110011",
		58 => "011001100100001110011",
		59 => "011001100100001110011",
		60 => "011000000100111010110",
		61 => "011000000100111010110",
		62 => "011000000100111010110",
		63 => "011001100100001010001",
		64 => "011001100100001010001",
		65 => "011001100100001010001",
		66 => "011001100100001110000",
		67 => "011001100100001110000",
		68 => "011001100100001110000",
		69 => "011001100100001010010",
		70 => "011001100100001010010",
		71 => "011001100100001010010",
		72 => "001000011100001010011",
		73 => "001000011100001010011",
		74 => "001000011100001010011",
		75 => "011001000100001010011",
		76 => "011001000100001010011",
		77 => "011001000100001010011",
		78 => "011000000100111010001",
		79 => "011000000100111010001",
		80 => "011000000100111010001",
		81 => "001000111101001010000",
		82 => "001000111101001010000",
		83 => "001000111101001010000",
		84 => "011000000101011010100",
		85 => "011000000101011010100",
		86 => "011000000101011010100",
		87 => "011010100100001010110",
		88 => "011010100100001010110",
		89 => "011010100100001010110",
		90 => "011000000110010011100",
		91 => "011000000110010011100",
		92 => "011000000110010011100",
		93 => "011101100100001011011",
		94 => "011101100100001011011",
		95 => "011101100100001011011",
		96 => "001001111100001010111",
		97 => "001001111100001010111",
		98 => "001001111100001010111",
		99 => "011000111100111010000",
		100 => "011000111100111010000",
		101 => "011000111100111010000",
		102 => "011000111100111010000",
		103 => "011000111100111010000",
		104 => "011000111100111010000",
		105 => "011001100100001110000",
		106 => "011001100100001110000",
		107 => "011001100100001110000",
		108 => "011000000101101010011",
		109 => "011000000101101010011",
		110 => "011000000101101010011",
		111 => "111000011101011010011",
		112 => "111000011101011010011",
		113 => "111000011101011010011",
		114 => "011000000101011010111",
		115 => "011000000101011010111",
		116 => "011000000101011010111",
		117 => "011000001100110110110",
		118 => "011000001100110110110",
		119 => "011000001100110110110",
		120 => "011011100100001010011",
		121 => "011011100100001010011",
		122 => "011011100100001010011",
		123 => "011000111100111010000",
		124 => "011000111100111010000",
		125 => "011000111100111010000",
		126 => "011000111100111010000",
		127 => "011000111100111010000",
		128 => "011000111100111010000",
		129 => "001000011100111010000",
		130 => "001000011100111010000",
		131 => "001000011100111010000",
		132 => "011000000101101010011",
		133 => "011000000101101010011",
		134 => "011000000101101010011",
		135 => "011000001101010010011",
		136 => "011000001101010010011",
		137 => "011000001101010010011",
		138 => "011000010100101011000",
		139 => "011000010100101011000",
		140 => "011000010100101011000",
		141 => "011000001100110110110",
		142 => "011000001100110110110",
		143 => "011000001100110110110",
		144 => "001001111100001010111",
		145 => "001001111100001010111",
		146 => "001001111100001010111",
		147 => "011000111100111010000",
		148 => "011000111100111010000",
		149 => "011000111100111010000",
		150 => "011000111100111010000",
		151 => "011000111100111010000",
		152 => "011000111100111010000",
		153 => "011001100100001110000",
		154 => "011001100100001110000",
		155 => "011001100100001110000",
		156 => "011000000101101010011",
		157 => "011000000101101010011",
		158 => "011000000101101010011",
		159 => "111000011101011010011",
		160 => "111000011101011010011",
		161 => "111000011101011010011",
		162 => "011000000101011010111",
		163 => "011000000101011010111",
		164 => "011000000101011010111",
		165 => "011000001100110110110",
		166 => "011000001100110110110",
		167 => "011000001100110110110",
		168 => "011011100100001010011",
		169 => "011011100100001010011",
		170 => "011011100100001010011",
		171 => "011000111100111010000",
		172 => "011000111100111010000",
		173 => "011000111100111010000",
		174 => "011000111100111010000",
		175 => "011000111100111010000",
		176 => "011000111100111010000",
		177 => "001000011100111010000",
		178 => "001000011100111010000",
		179 => "001000011100111010000",
		180 => "011000000101101010011",
		181 => "011000000101101010011",
		182 => "011000000101101010011",
		183 => "011000001101010010011",
		184 => "011000001101010010011",
		185 => "011000001101010010011",
		186 => "011000010100101011000",
		187 => "011000010100101011000",
		188 => "011000010100101011000",
		189 => "011000001100110110110",
		190 => "011000001100110110110",
		191 => "011000001100110110110",
		192 => "001001100101101110000",
		193 => "001001100101101110000",
		194 => "001001100101101110000",
		195 => "011000001100101010110",
		196 => "011000001100101010110",
		197 => "011000001100101010110",
		198 => "011000000100111010001",
		199 => "011000000100111010001",
		200 => "011000000100111010001",
		201 => "001001111110001010000",
		202 => "001001111110001010000",
		203 => "001001111110001010000",
		204 => "001000010100111010110",
		205 => "001000010100111010110",
		206 => "001000010100111010110",
		207 => "001000111100011110011",
		208 => "001000111100011110011",
		209 => "001000111100011110011",
		210 => "011000000100111010001",
		211 => "011000000100111010001",
		212 => "011000000100111010001",
		213 => "001001111110001010000",
		214 => "001001111110001010000",
		215 => "001001111110001010000",
		216 => "001001100101101110000",
		217 => "001001100101101110000",
		218 => "001001100101101110000",
		219 => "011000001100101010110",
		220 => "011000001100101010110",
		221 => "011000001100101010110",
		222 => "011000000100111010001",
		223 => "011000000100111010001",
		224 => "011000000100111010001",
		225 => "001001111110001010000",
		226 => "001001111110001010000",
		227 => "001001111110001010000",
		228 => "001000010100111010110",
		229 => "001000010100111010110",
		230 => "001000010100111010110",
		231 => "001000111100011110011",
		232 => "001000111100011110011",
		233 => "001000111100011110011",
		234 => "011000000100111010001",
		235 => "011000000100111010001",
		236 => "011000000100111010001",
		237 => "001001111110001010000",
		238 => "001001111110001010000",
		239 => "001001111110001010000",
		240 => "001001100101101110000",
		241 => "001001100101101110000",
		242 => "001001100101101110000",
		243 => "011000001100101010110",
		244 => "011000001100101010110",
		245 => "011000001100101010110",
		246 => "011000000100111010001",
		247 => "011000000100111010001",
		248 => "011000000100111010001",
		249 => "001001111110001010000",
		250 => "001001111110001010000",
		251 => "001001111110001010000",
		252 => "001000010100111010110",
		253 => "001000010100111010110",
		254 => "001000010100111010110",
		255 => "001000111100011110011",
		256 => "001000111100011110011",
		257 => "001000111100011110011",
		258 => "011000000100111010001",
		259 => "011000000100111010001",
		260 => "011000000100111010001",
		261 => "001001111110001010000",
		262 => "001001111110001010000",
		263 => "001001111110001010000",
		264 => "001001100101101110000",
		265 => "001001100101101110000",
		266 => "001001100101101110000",
		267 => "011000001100101010110",
		268 => "011000001100101010110",
		269 => "011000001100101010110",
		270 => "011000000100111010001",
		271 => "011000000100111010001",
		272 => "011000000100111010001",
		273 => "001001111110001010000",
		274 => "001001111110001010000",
		275 => "001001111110001010000",
		276 => "001000010100111010110",
		277 => "001000010100111010110",
		278 => "001000010100111010110",
		279 => "001000111100011110011",
		280 => "001000111100011110011",
		281 => "001000111100011110011",
		282 => "011000000100111010001",
		283 => "011000000100111010001",
		284 => "011000000100111010001",
		285 => "001001111110001010000",
		286 => "001001111110001010000",
		287 => "001001111110001010000",
		288 => "001011011100001010111",
		289 => "001011011100001010111",
		290 => "001011011100001010111",
		291 => "011000001110100010101",
		292 => "011000001110100010101",
		293 => "011000001110100010101",
		294 => "011000111100111010000",
		295 => "011000111100111010000",
		296 => "011000111100111010000",
		297 => "011000001110100010101",
		298 => "011000001110100010101",
		299 => "011000001110100010101",
		300 => "001011011100001010111",
		301 => "001011011100001010111",
		302 => "001011011100001010111",
		303 => "011000001110100010101",
		304 => "011000001110100010101",
		305 => "011000001110100010101",
		306 => "011000111100111010000",
		307 => "011000111100111010000",
		308 => "011000111100111010000",
		309 => "011000001110100010101",
		310 => "011000001110100010101",
		311 => "011000001110100010101",
		312 => "001011011100001010111",
		313 => "001011011100001010111",
		314 => "001011011100001010111",
		315 => "011000001110100010101",
		316 => "011000001110100010101",
		317 => "011000001110100010101",
		318 => "011000111100111010000",
		319 => "011000111100111010000",
		320 => "011000111100111010000",
		321 => "011000001110100010101",
		322 => "011000001110100010101",
		323 => "011000001110100010101",
		324 => "001011011100001010111",
		325 => "001011011100001010111",
		326 => "001011011100001010111",
		327 => "011000001110100010101",
		328 => "011000001110100010101",
		329 => "011000001110100010101",
		330 => "011000111100111010000",
		331 => "011000111100111010000",
		332 => "011000111100111010000",
		333 => "011000001110100010101",
		334 => "011000001110100010101",
		335 => "011000001110100010101",
		336 => "001011011100001010111",
		337 => "001011011100001010111",
		338 => "001011011100001010111",
		339 => "011000001110100010101",
		340 => "011000001110100010101",
		341 => "011000001110100010101",
		342 => "011000111100111010000",
		343 => "011000111100111010000",
		344 => "011000111100111010000",
		345 => "011000001110100010101",
		346 => "011000001110100010101",
		347 => "011000001110100010101",
		348 => "001011011100001010111",
		349 => "001011011100001010111",
		350 => "001011011100001010111",
		351 => "011000001110100010101",
		352 => "011000001110100010101",
		353 => "011000001110100010101",
		354 => "011000111100111010000",
		355 => "011000111100111010000",
		356 => "011000111100111010000",
		357 => "011000001110100010101",
		358 => "011000001110100010101",
		359 => "011000001110100010101",
		360 => "001011011100001010111",
		361 => "001011011100001010111",
		362 => "001011011100001010111",
		363 => "011000001110100010101",
		364 => "011000001110100010101",
		365 => "011000001110100010101",
		366 => "011000111100111010000",
		367 => "011000111100111010000",
		368 => "011000111100111010000",
		369 => "011000001110100010101",
		370 => "011000001110100010101",
		371 => "011000001110100010101",
		372 => "001011011100001010111",
		373 => "001011011100001010111",
		374 => "001011011100001010111",
		375 => "011000001110100010101",
		376 => "011000001110100010101",
		377 => "011000001110100010101",
		378 => "011000111100111010000",
		379 => "011000111100111010000",
		380 => "011000111100111010000",
		381 => "011000001110100010101",
		382 => "011000001110100010101",
		383 => "011000001110100010101",
		384 => "011001011100001010100",
		385 => "011001011100001010100",
		386 => "011001011100001010100",
		387 => "011010000100001110010",
		388 => "011010000100001110010",
		389 => "011010000100001110010",
		390 => "011001011100001010100",
		391 => "011001011100001010100",
		392 => "011001011100001010100",
		393 => "011010000100001110010",
		394 => "011010000100001110010",
		395 => "011010000100001110010",
		396 => "011001011100001010100",
		397 => "011001011100001010100",
		398 => "011001011100001010100",
		399 => "011010000100001110010",
		400 => "011010000100001110010",
		401 => "011010000100001110010",
		402 => "011001011100001010100",
		403 => "011001011100001010100",
		404 => "011001011100001010100",
		405 => "011010000100001110010",
		406 => "011010000100001110010",
		407 => "011010000100001110010",
		408 => "011001011100001010100",
		409 => "011001011100001010100",
		410 => "011001011100001010100",
		411 => "011010000100001110010",
		412 => "011010000100001110010",
		413 => "011010000100001110010",
		414 => "011001011100001010100",
		415 => "011001011100001010100",
		416 => "011001011100001010100",
		417 => "011010000100001110010",
		418 => "011010000100001110010",
		419 => "011010000100001110010",
		420 => "011001011100001010100",
		421 => "011001011100001010100",
		422 => "011001011100001010100",
		423 => "011010000100001110010",
		424 => "011010000100001110010",
		425 => "011010000100001110010",
		426 => "011001011100001010100",
		427 => "011001011100001010100",
		428 => "011001011100001010100",
		429 => "011010000100001110010",
		430 => "011010000100001110010",
		431 => "011010000100001110010",
		432 => "011001011100001010100",
		433 => "011001011100001010100",
		434 => "011001011100001010100",
		435 => "011010000100001110010",
		436 => "011010000100001110010",
		437 => "011010000100001110010",
		438 => "011001011100001010100",
		439 => "011001011100001010100",
		440 => "011001011100001010100",
		441 => "011010000100001110010",
		442 => "011010000100001110010",
		443 => "011010000100001110010",
		444 => "011001011100001010100",
		445 => "011001011100001010100",
		446 => "011001011100001010100",
		447 => "011010000100001110010",
		448 => "011010000100001110010",
		449 => "011010000100001110010",
		450 => "011001011100001010100",
		451 => "011001011100001010100",
		452 => "011001011100001010100",
		453 => "011010000100001110010",
		454 => "011010000100001110010",
		455 => "011010000100001110010",
		456 => "011001011100001010100",
		457 => "011001011100001010100",
		458 => "011001011100001010100",
		459 => "011010000100001110010",
		460 => "011010000100001110010",
		461 => "011010000100001110010",
		462 => "011001011100001010100",
		463 => "011001011100001010100",
		464 => "011001011100001010100",
		465 => "011010000100001110010",
		466 => "011010000100001110010",
		467 => "011010000100001110010",
		468 => "011001011100001010100",
		469 => "011001011100001010100",
		470 => "011001011100001010100",
		471 => "011010000100001110010",
		472 => "011010000100001110010",
		473 => "011010000100001110010",
		474 => "011001011100001010100",
		475 => "011001011100001010100",
		476 => "011001011100001010100",
		477 => "011010000100001110010",
		478 => "011010000100001110010",
		479 => "011010000100001110010",
		480 => "011000001101100010011",
		481 => "011000001101100010011",
		482 => "011000001101100010011",
		483 => "011000001101100010011",
		484 => "011000001101100010011",
		485 => "011000001101100010011",
		486 => "011000001101100010011",
		487 => "011000001101100010011",
		488 => "011000001101100010011",
		489 => "011000001101100010011",
		490 => "011000001101100010011",
		491 => "011000001101100010011",
		492 => "011000001101100010011",
		493 => "011000001101100010011",
		494 => "011000001101100010011",
		495 => "011000001101100010011",
		496 => "011000001101100010011",
		497 => "011000001101100010011",
		498 => "011000001101100010011",
		499 => "011000001101100010011",
		500 => "011000001101100010011",
		501 => "011000001101100010011",
		502 => "011000001101100010011",
		503 => "011000001101100010011",
		504 => "011000001101100010011",
		505 => "011000001101100010011",
		506 => "011000001101100010011",
		507 => "011000001101100010011",
		508 => "011000001101100010011",
		509 => "011000001101100010011",
		510 => "011000001101100010011",
		511 => "011000001101100010011",
		512 => "011000001101100010011",
		513 => "011000001101100010011",
		514 => "011000001101100010011",
		515 => "011000001101100010011",
		516 => "011000001101100010011",
		517 => "011000001101100010011",
		518 => "011000001101100010011",
		519 => "011000001101100010011",
		520 => "011000001101100010011",
		521 => "011000001101100010011",
		522 => "011000001101100010011",
		523 => "011000001101100010011",
		524 => "011000001101100010011",
		525 => "011000001101100010011",
		526 => "011000001101100010011",
		527 => "011000001101100010011",
		528 => "011000001101100010011",
		529 => "011000001101100010011",
		530 => "011000001101100010011",
		531 => "011000001101100010011",
		532 => "011000001101100010011",
		533 => "011000001101100010011",
		534 => "011000001101100010011",
		535 => "011000001101100010011",
		536 => "011000001101100010011",
		537 => "011000001101100010011",
		538 => "011000001101100010011",
		539 => "011000001101100010011",
		540 => "011000001101100010011",
		541 => "011000001101100010011",
		542 => "011000001101100010011",
		543 => "011000001101100010011",
		544 => "011000001101100010011",
		545 => "011000001101100010011",
		546 => "011000001101100010011",
		547 => "011000001101100010011",
		548 => "011000001101100010011",
		549 => "011000001101100010011",
		550 => "011000001101100010011",
		551 => "011000001101100010011",
		552 => "011000001101100010011",
		553 => "011000001101100010011",
		554 => "011000001101100010011",
		555 => "011000001101100010011",
		556 => "011000001101100010011",
		557 => "011000001101100010011",
		558 => "011000001101100010011",
		559 => "011000001101100010011",
		560 => "011000001101100010011",
		561 => "011000001101100010011",
		562 => "011000001101100010011",
		563 => "011000001101100010011",
		564 => "011000001101100010011",
		565 => "011000001101100010011",
		566 => "011000001101100010011",
		567 => "011000001101100010011",
		568 => "011000001101100010011",
		569 => "011000001101100010011",
		570 => "011000001101100010011",
		571 => "011000001101100010011",
		572 => "011000001101100010011",
		573 => "011000001101100010011",
		574 => "011000001101100010011",
		575 => "011000001101100010011",
		576 => "011001100100001110001",
		577 => "011001100100001110001",
		578 => "011001100100001110001",
		579 => "011001100100001110001",
		580 => "011001100100001110001",
		581 => "011001100100001110001",
		582 => "011001100100001110001",
		583 => "011001100100001110001",
		584 => "011001100100001110001",
		585 => "011001100100001110001",
		586 => "011001100100001110001",
		587 => "011001100100001110001",
		588 => "011001100100001110001",
		589 => "011001100100001110001",
		590 => "011001100100001110001",
		591 => "011001100100001110001",
		592 => "011001100100001110001",
		593 => "011001100100001110001",
		594 => "011001100100001110001",
		595 => "011001100100001110001",
		596 => "011001100100001110001",
		597 => "011001100100001110001",
		598 => "011001100100001110001",
		599 => "011001100100001110001",
		600 => "011001100100001110001",
		601 => "011001100100001110001",
		602 => "011001100100001110001",
		603 => "011001100100001110001",
		604 => "011001100100001110001",
		605 => "011001100100001110001",
		606 => "011001100100001110001",
		607 => "011001100100001110001",
		608 => "011001100100001110001",
		609 => "011001100100001110001",
		610 => "011001100100001110001",
		611 => "011001100100001110001",
		612 => "011001100100001110001",
		613 => "011001100100001110001",
		614 => "011001100100001110001",
		615 => "011001100100001110001",
		616 => "011001100100001110001",
		617 => "011001100100001110001",
		618 => "011001100100001110001",
		619 => "011001100100001110001",
		620 => "011001100100001110001",
		621 => "011001100100001110001",
		622 => "011001100100001110001",
		623 => "011001100100001110001",
		624 => "011001100100001110001",
		625 => "011001100100001110001",
		626 => "011001100100001110001",
		627 => "011001100100001110001",
		628 => "011001100100001110001",
		629 => "011001100100001110001",
		630 => "011001100100001110001",
		631 => "011001100100001110001",
		632 => "011001100100001110001",
		633 => "011001100100001110001",
		634 => "011001100100001110001",
		635 => "011001100100001110001",
		636 => "011001100100001110001",
		637 => "011001100100001110001",
		638 => "011001100100001110001",
		639 => "011001100100001110001",
		640 => "011001100100001110001",
		641 => "011001100100001110001",
		642 => "011001100100001110001",
		643 => "011001100100001110001",
		644 => "011001100100001110001",
		645 => "011001100100001110001",
		646 => "011001100100001110001",
		647 => "011001100100001110001",
		648 => "011001100100001110001",
		649 => "011001100100001110001",
		650 => "011001100100001110001",
		651 => "011001100100001110001",
		652 => "011001100100001110001",
		653 => "011001100100001110001",
		654 => "011001100100001110001",
		655 => "011001100100001110001",
		656 => "011001100100001110001",
		657 => "011001100100001110001",
		658 => "011001100100001110001",
		659 => "011001100100001110001",
		660 => "011001100100001110001",
		661 => "011001100100001110001",
		662 => "011001100100001110001",
		663 => "011001100100001110001",
		664 => "011001100100001110001",
		665 => "011001100100001110001",
		666 => "011001100100001110001",
		667 => "011001100100001110001",
		668 => "011001100100001110001",
		669 => "011001100100001110001",
		670 => "011001100100001110001",
		671 => "011001100100001110001",
		672 => "011000101100100010101",
		673 => "011000101100100010101",
		674 => "011000101100100010101",
		675 => "011000101100100010101",
		676 => "011000101100100010101",
		677 => "011000101100100010101",
		678 => "011000101100100010101",
		679 => "011000101100100010101",
		680 => "011000101100100010101",
		681 => "011000101100100010101",
		682 => "011000101100100010101",
		683 => "011000101100100010101",
		684 => "011000101100100010101",
		685 => "011000101100100010101",
		686 => "011000101100100010101",
		687 => "011000101100100010101",
		688 => "011000101100100010101",
		689 => "011000101100100010101",
		690 => "011000101100100010101",
		691 => "011000101100100010101",
		692 => "011000101100100010101",
		693 => "011000101100100010101",
		694 => "011000101100100010101",
		695 => "011000101100100010101",
		696 => "011000101100100010101",
		697 => "011000101100100010101",
		698 => "011000101100100010101",
		699 => "011000101100100010101",
		700 => "011000101100100010101",
		701 => "011000101100100010101",
		702 => "011000101100100010101",
		703 => "011000101100100010101",
		704 => "011000101100100010101",
		705 => "011000101100100010101",
		706 => "011000101100100010101",
		707 => "011000101100100010101",
		708 => "011000101100100010101",
		709 => "011000101100100010101",
		710 => "011000101100100010101",
		711 => "011000101100100010101",
		712 => "011000101100100010101",
		713 => "011000101100100010101",
		714 => "011000101100100010101",
		715 => "011000101100100010101",
		716 => "011000101100100010101",
		717 => "011000101100100010101",
		718 => "011000101100100010101",
		719 => "011000101100100010101",
		720 => "011000101100100010101",
		721 => "011000101100100010101",
		722 => "011000101100100010101",
		723 => "011000101100100010101",
		724 => "011000101100100010101",
		725 => "011000101100100010101",
		726 => "011000101100100010101",
		727 => "011000101100100010101",
		728 => "011000101100100010101",
		729 => "011000101100100010101",
		730 => "011000101100100010101",
		731 => "011000101100100010101",
		732 => "011000101100100010101",
		733 => "011000101100100010101",
		734 => "011000101100100010101",
		735 => "011000101100100010101",
		736 => "011000101100100010101",
		737 => "011000101100100010101",
		738 => "011000101100100010101",
		739 => "011000101100100010101",
		740 => "011000101100100010101",
		741 => "011000101100100010101",
		742 => "011000101100100010101",
		743 => "011000101100100010101",
		744 => "011000101100100010101",
		745 => "011000101100100010101",
		746 => "011000101100100010101",
		747 => "011000101100100010101",
		748 => "011000101100100010101",
		749 => "011000101100100010101",
		750 => "011000101100100010101",
		751 => "011000101100100010101",
		752 => "011000101100100010101",
		753 => "011000101100100010101",
		754 => "011000101100100010101",
		755 => "011000101100100010101",
		756 => "011000101100100010101",
		757 => "011000101100100010101",
		758 => "011000101100100010101",
		759 => "011000101100100010101",
		760 => "011000101100100010101",
		761 => "011000101100100010101",
		762 => "011000101100100010101",
		763 => "011000101100100010101",
		764 => "011000101100100010101",
		765 => "011000101100100010101",
		766 => "011000101100100010101",
		767 => "011000101100100010101",
		768 => "011000101100100110010",
		769 => "011000101100100110010",
		770 => "011000101100100110010",
		771 => "011000101100100110010",
		772 => "011000101100100110010",
		773 => "011000101100100110010",
		774 => "011000101100100110010",
		775 => "011000101100100110010",
		776 => "011000101100100110010",
		777 => "011000101100100110010",
		778 => "011000101100100110010",
		779 => "011000101100100110010",
		780 => "011000101100100110010",
		781 => "011000101100100110010",
		782 => "011000101100100110010",
		783 => "011000101100100110010",
		784 => "011000101100100110010",
		785 => "011000101100100110010",
		786 => "011000101100100110010",
		787 => "011000101100100110010",
		788 => "011000101100100110010",
		789 => "011000101100100110010",
		790 => "011000101100100110010",
		791 => "011000101100100110010",
		792 => "011000101100100110010",
		793 => "011000101100100110010",
		794 => "011000101100100110010",
		795 => "011000101100100110010",
		796 => "011000101100100110010",
		797 => "011000101100100110010",
		798 => "011000101100100110010",
		799 => "011000101100100110010",
		800 => "011000101100100110010",
		801 => "011000101100100110010",
		802 => "011000101100100110010",
		803 => "011000101100100110010",
		804 => "011000101100100110010",
		805 => "011000101100100110010",
		806 => "011000101100100110010",
		807 => "011000101100100110010",
		808 => "011000101100100110010",
		809 => "011000101100100110010",
		810 => "011000101100100110010",
		811 => "011000101100100110010",
		812 => "011000101100100110010",
		813 => "011000101100100110010",
		814 => "011000101100100110010",
		815 => "011000101100100110010",
		816 => "011000101100100110010",
		817 => "011000101100100110010",
		818 => "011000101100100110010",
		819 => "011000101100100110010",
		820 => "011000101100100110010",
		821 => "011000101100100110010",
		822 => "011000101100100110010",
		823 => "011000101100100110010",
		824 => "011000101100100110010",
		825 => "011000101100100110010",
		826 => "011000101100100110010",
		827 => "011000101100100110010",
		828 => "011000101100100110010",
		829 => "011000101100100110010",
		830 => "011000101100100110010",
		831 => "011000101100100110010",
		832 => "011000101100100110010",
		833 => "011000101100100110010",
		834 => "011000101100100110010",
		835 => "011000101100100110010",
		836 => "011000101100100110010",
		837 => "011000101100100110010",
		838 => "011000101100100110010",
		839 => "011000101100100110010",
		840 => "011000101100100110010",
		841 => "011000101100100110010",
		842 => "011000101100100110010",
		843 => "011000101100100110010",
		844 => "011000101100100110010",
		845 => "011000101100100110010",
		846 => "011000101100100110010",
		847 => "011000101100100110010",
		848 => "011000101100100110010",
		849 => "011000101100100110010",
		850 => "011000101100100110010",
		851 => "011000101100100110010",
		852 => "011000101100100110010",
		853 => "011000101100100110010",
		854 => "011000101100100110010",
		855 => "011000101100100110010",
		856 => "011000101100100110010",
		857 => "011000101100100110010",
		858 => "011000101100100110010",
		859 => "011000101100100110010",
		860 => "011000101100100110010",
		861 => "011000101100100110010",
		862 => "011000101100100110010",
		863 => "011000101100100110010");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;