LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.MainPackage.all;

ENTITY DisplayMod IS
	PORT(Clock: IN STD_LOGIC;
		  reset: IN STD_LOGIC;
		  CurrentState: IN StateFFT;
		  SF_D : OUT STD_LOGIC_VECTOR(3 downto 0);
		  LCD_E: OUT STD_LOGIC;
		  LCD_RS: OUT STD_LOGIC;
		  LCD_RW: OUT STD_LOGIC);
END DisplayMod;

ARCHITECTURE Logica OF DisplayMod IS
	
	CONSTANT ResetDisplay : INFO :=        ("10100000","01000110","01000110","01010100","10100000","01010010","01000001","01000100","01001001","01011000","00101101","00110010","10100000","00111000","01010000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000");
	CONSTANT IdleDisplay : INFO :=         ("10100000","01000110","01000110","01010100","10100000","01010010","01000001","01000100","01001001","01011000","00101101","00110010","10100000","00111000","01010000","10100000","10100000","01000101","01101101","10100000","01000101","01110011","01110000","01100101","01110010","01100001","10100000","10100000","10100000","10100000","10100000","10100000");
	CONSTANT ReceiveDataDisplay : INFO :=  ("10100000","01000110","01000110","01010100","10100000","01010010","01000001","01000100","01001001","01011000","00101101","00110010","10100000","00111000","01010000","10100000","10100000","01010010","01100101","01100011","01100101","01100011","01100101","01101110","01100100","01101111","10100000","01000100","01100001","01100100","01101111","01110011");
	CONSTANT ProcessDataDisplay : INFO :=  ("10100000","01000110","01000110","01010100","10100000","01010010","01000001","01000100","01001001","01011000","00101101","00110010","10100000","00111000","01010000","10100000","10100000","01000011","01100001","01101100","01100011","01110101","01101100","01100001","01101110","01100100","01101111","10100000","01000110","01000110","01010100","10100000");
	CONSTANT TransmitDataDisplay : INFO := ("10100000","01000110","01000110","01010100","10100000","01010010","01000001","01000100","01001001","01011000","00101101","00110010","10100000","00111000","01010000","10100000","10100000","01000101","01101110","01110110","01101001","01100001","01101110","01100100","01101111","10100000","01000100","01100001","01100100","01101111","01110011","10100000");
	SIGNAL RstDisplay : STD_LOGIC := '0';
	SIGNAL DATA: INFO := ("10100000","01000110","01000110","01010100","10100000","01010010","01000001","01000100","01001001","01011000","00101101","00110010","10100000","00111000","01010000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000","10100000");
	                   --(  BLANK        F          F          T        BLANK        R           A         D          I          X         -          2         BLANK        8           P       BLANK     BLANK        BLANK     BLANK       BLANK     BLANK        BLANK     BLANK     BLANK     BLANK        BLANK     BLANK       BLANK     BLANK        BLANK     BLANK     BLANK 
							 --(     1         2          3          4          5          6           7         8          9          10        11         12           13       14          15         16         17         18         19         20         21         22         23        24           25       26         27          28         29       30          31          32  
	
	BEGIN
	
	---------------------------------------------------------------
	--               Dispositivo de Print na tela                --
	---------------------------------------------------------------	
	Display: DisplayLCD PORT MAP(Clock,reset, RstDisplay, DATA, SF_D,LCD_E,LCD_RS,LCD_RW);	
	
	
	---------------------------------------------------------------
	--                       Sele��o de Data                     --
	---------------------------------------------------------------
	DATA <=  ResetDisplay        WHEN CurrentState = ResetFFT     ELSE
			   IdleDisplay         WHEN CurrentState = Idle         ELSE
			   ReceiveDataDisplay  WHEN CurrentState = ReceiveData  ELSE
			   ProcessDataDisplay  WHEN CurrentState = ProcessData  ELSE
			   TransmitDataDisplay WHEN CurrentState = TransmitData;
				
	---------------------------------------------------------------
	--               Dispositivo de Print na tela                --
	---------------------------------------------------------------
	Trigger : PROCESS(reset, Clock)
	
		VARIABLE Actual: StateFFT ;
		VARIABLE Before: StateFFT ;
	
	BEGIN
	
		IF(reset = '1') THEN
			RstDisplay <= '0';
		
		ELSIF(clock = '1' AND clock'EVENT) THEN
			Actual := CurrentState;
			IF(Actual /= Before) THEN
				Before := CurrentState;
				RstDisplay <= '1';
				
			ELSE
				RstDisplay <= '0';
				
			END IF;
			
		END IF;
	
	END PROCESS;

END Logica;
