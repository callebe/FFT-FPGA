library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT2 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT2;

architecture Behavioral of ROMFFT2 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 3 
	constant ROM_tb : ROM := (
		0 => "011011000110111010000",
		1 => "011011000110111010000",
		2 => "011011000110111010000",
		3 => "011000000101111010110",
		4 => "011000000101111010110",
		5 => "011000000101111010110",
		6 => "011010100100001110101",
		7 => "011010100100001110101",
		8 => "011010100100001110101",
		9 => "011010100100001010100",
		10 => "011010100100001010100",
		11 => "011010100100001010100",
		12 => "011001011100111010000",
		13 => "011001011100111010000",
		14 => "011001011100111010000",
		15 => "001001011100001010101",
		16 => "001001011100001010101",
		17 => "001001011100001010101",
		18 => "001000111100001110110",
		19 => "001000111100001110110",
		20 => "001000111100001110110",
		21 => "001010111100001110010",
		22 => "001010111100001110010",
		23 => "001010111100001110010",
		24 => "011001100100001110000",
		25 => "011001100100001110000",
		26 => "011001100100001110000",
		27 => "011000101100111010001",
		28 => "011000101100111010001",
		29 => "011000101100111010001",
		30 => "011000010100011010011",
		31 => "011000010100011010011",
		32 => "011000010100011010011",
		33 => "011000000100111010110",
		34 => "011000000100111010110",
		35 => "011000000100111010110",
		36 => "011000001100101010001",
		37 => "011000001100101010001",
		38 => "011000001100101010001",
		39 => "011000000101011010011",
		40 => "011000000101011010011",
		41 => "011000000101011010011",
		42 => "011000000101111010100",
		43 => "011000000101111010100",
		44 => "011000000101111010100",
		45 => "011010111100001011001",
		46 => "011010111100001011001",
		47 => "011010111100001011001",
		48 => "011101100101101110000",
		49 => "011101100101101110000",
		50 => "011101100101101110000",
		51 => "011000000101111010110",
		52 => "011000000101111010110",
		53 => "011000000101111010110",
		54 => "011010100100001110101",
		55 => "011010100100001110101",
		56 => "011010100100001110101",
		57 => "011010100100001010100",
		58 => "011010100100001010100",
		59 => "011010100100001010100",
		60 => "011001011100111010000",
		61 => "011001011100111010000",
		62 => "011001011100111010000",
		63 => "011010100100001010010",
		64 => "011010100100001010010",
		65 => "011010100100001010010",
		66 => "001000000101101010001",
		67 => "001000000101101010001",
		68 => "001000000101101010001",
		69 => "001000000100101010101",
		70 => "001000000100101010101",
		71 => "001000000100101010101",
		72 => "001000011100111010000",
		73 => "001000011100111010000",
		74 => "001000011100111010000",
		75 => "011000101100111010001",
		76 => "011000101100111010001",
		77 => "011000101100111010001",
		78 => "011000010100011010011",
		79 => "011000010100011010011",
		80 => "011000010100011010011",
		81 => "011000000100111010110",
		82 => "011000000100111010110",
		83 => "011000000100111010110",
		84 => "001000000100101110001",
		85 => "001000000100101110001",
		86 => "001000000100101110001",
		87 => "011010100100001110011",
		88 => "011010100100001110011",
		89 => "011010100100001110011",
		90 => "001010011101111010000",
		91 => "001010011101111010000",
		92 => "001010011101111010000",
		93 => "011100100100001110101",
		94 => "011100100100001110101",
		95 => "011100100100001110101",
		96 => "011000000110111110101",
		97 => "011000000110111110101",
		98 => "011000000110111110101",
		99 => "011010100100001010010",
		100 => "011010100100001010010",
		101 => "011010100100001010010",
		102 => "001000111100001110011",
		103 => "001000111100001110011",
		104 => "001000111100001110011",
		105 => "011001111100011110010",
		106 => "011001111100011110010",
		107 => "011001111100011110010",
		108 => "011001100100001110000",
		109 => "011001100100001110000",
		110 => "011001100100001110000",
		111 => "011000000101001010010",
		112 => "011000000101001010010",
		113 => "011000000101001010010",
		114 => "011010100100001110010",
		115 => "011010100100001110010",
		116 => "011010100100001110010",
		117 => "011000000101111010100",
		118 => "011000000101111010100",
		119 => "011000000101111010100",
		120 => "001010111100001011011",
		121 => "001010111100001011011",
		122 => "001010111100001011011",
		123 => "001001011100001010101",
		124 => "001001011100001010101",
		125 => "001001011100001010101",
		126 => "001000111100001110011",
		127 => "001000111100001110011",
		128 => "001000111100001110011",
		129 => "011001000100001110011",
		130 => "011001000100001110011",
		131 => "011001000100001110011",
		132 => "001000011100111010000",
		133 => "001000011100111010000",
		134 => "001000011100111010000",
		135 => "011000000101001010010",
		136 => "011000000101001010010",
		137 => "011000000101001010010",
		138 => "011000000101011010010",
		139 => "011000000101011010010",
		140 => "011000000101011010010",
		141 => "011011100100001110100",
		142 => "011011100100001110100",
		143 => "011011100100001110100",
		144 => "011000000110111110101",
		145 => "011000000110111110101",
		146 => "011000000110111110101",
		147 => "011010100100001010010",
		148 => "011010100100001010010",
		149 => "011010100100001010010",
		150 => "001000111100001110011",
		151 => "001000111100001110011",
		152 => "001000111100001110011",
		153 => "011001111100011110010",
		154 => "011001111100011110010",
		155 => "011001111100011110010",
		156 => "011001100100001110000",
		157 => "011001100100001110000",
		158 => "011001100100001110000",
		159 => "011000000101001010010",
		160 => "011000000101001010010",
		161 => "011000000101001010010",
		162 => "011010100100001110010",
		163 => "011010100100001110010",
		164 => "011010100100001110010",
		165 => "011000000101111010100",
		166 => "011000000101111010100",
		167 => "011000000101111010100",
		168 => "001010111100001011011",
		169 => "001010111100001011011",
		170 => "001010111100001011011",
		171 => "001001011100001010101",
		172 => "001001011100001010101",
		173 => "001001011100001010101",
		174 => "001000111100001110011",
		175 => "001000111100001110011",
		176 => "001000111100001110011",
		177 => "011001000100001110011",
		178 => "011001000100001110011",
		179 => "011001000100001110011",
		180 => "001000011100111010000",
		181 => "001000011100111010000",
		182 => "001000011100111010000",
		183 => "011000000101001010010",
		184 => "011000000101001010010",
		185 => "011000000101001010010",
		186 => "011000000101011010010",
		187 => "011000000101011010010",
		188 => "011000000101011010010",
		189 => "011011100100001110100",
		190 => "011011100100001110100",
		191 => "011011100100001110100",
		192 => "011000000110011110100",
		193 => "011000000110011110100",
		194 => "011000000110011110100",
		195 => "011000000100111010110",
		196 => "011000000100111010110",
		197 => "011000000100111010110",
		198 => "011001011100001010011",
		199 => "011001011100001010011",
		200 => "011001011100001010011",
		201 => "011000000101011010011",
		202 => "011000000101011010011",
		203 => "011000000101011010011",
		204 => "001010011100001011001",
		205 => "001010011100001011001",
		206 => "001010011100001011001",
		207 => "011000001101110010011",
		208 => "011000001101110010011",
		209 => "011000001101110010011",
		210 => "011001100100001110010",
		211 => "011001100100001110010",
		212 => "011001100100001110010",
		213 => "011010100100001110011",
		214 => "011010100100001110011",
		215 => "011010100100001110011",
		216 => "011000000110011110100",
		217 => "011000000110011110100",
		218 => "011000000110011110100",
		219 => "011000000100111010110",
		220 => "011000000100111010110",
		221 => "011000000100111010110",
		222 => "011001011100001010011",
		223 => "011001011100001010011",
		224 => "011001011100001010011",
		225 => "011000000101011010011",
		226 => "011000000101011010011",
		227 => "011000000101011010011",
		228 => "001010011100001011001",
		229 => "001010011100001011001",
		230 => "001010011100001011001",
		231 => "011000001101110010011",
		232 => "011000001101110010011",
		233 => "011000001101110010011",
		234 => "011001100100001110010",
		235 => "011001100100001110010",
		236 => "011001100100001110010",
		237 => "011010100100001110011",
		238 => "011010100100001110011",
		239 => "011010100100001110011",
		240 => "011000000110011110100",
		241 => "011000000110011110100",
		242 => "011000000110011110100",
		243 => "011000000100111010110",
		244 => "011000000100111010110",
		245 => "011000000100111010110",
		246 => "011001011100001010011",
		247 => "011001011100001010011",
		248 => "011001011100001010011",
		249 => "011000000101011010011",
		250 => "011000000101011010011",
		251 => "011000000101011010011",
		252 => "001010011100001011001",
		253 => "001010011100001011001",
		254 => "001010011100001011001",
		255 => "011000001101110010011",
		256 => "011000001101110010011",
		257 => "011000001101110010011",
		258 => "011001100100001110010",
		259 => "011001100100001110010",
		260 => "011001100100001110010",
		261 => "011010100100001110011",
		262 => "011010100100001110011",
		263 => "011010100100001110011",
		264 => "011000000110011110100",
		265 => "011000000110011110100",
		266 => "011000000110011110100",
		267 => "011000000100111010110",
		268 => "011000000100111010110",
		269 => "011000000100111010110",
		270 => "011001011100001010011",
		271 => "011001011100001010011",
		272 => "011001011100001010011",
		273 => "011000000101011010011",
		274 => "011000000101011010011",
		275 => "011000000101011010011",
		276 => "001010011100001011001",
		277 => "001010011100001011001",
		278 => "001010011100001011001",
		279 => "011000001101110010011",
		280 => "011000001101110010011",
		281 => "011000001101110010011",
		282 => "011001100100001110010",
		283 => "011001100100001110010",
		284 => "011001100100001110010",
		285 => "011010100100001110011",
		286 => "011010100100001110011",
		287 => "011010100100001110011",
		288 => "011000000101111110011",
		289 => "011000000101111110011",
		290 => "011000000101111110011",
		291 => "011000101100111010001",
		292 => "011000101100111010001",
		293 => "011000101100111010001",
		294 => "001001111100001010111",
		295 => "001001111100001010111",
		296 => "001001111100001010111",
		297 => "001000000100101110110",
		298 => "001000000100101110110",
		299 => "001000000100101110110",
		300 => "011000000101111110011",
		301 => "011000000101111110011",
		302 => "011000000101111110011",
		303 => "011000101100111010001",
		304 => "011000101100111010001",
		305 => "011000101100111010001",
		306 => "001001111100001010111",
		307 => "001001111100001010111",
		308 => "001001111100001010111",
		309 => "001000000100101110110",
		310 => "001000000100101110110",
		311 => "001000000100101110110",
		312 => "011000000101111110011",
		313 => "011000000101111110011",
		314 => "011000000101111110011",
		315 => "011000101100111010001",
		316 => "011000101100111010001",
		317 => "011000101100111010001",
		318 => "001001111100001010111",
		319 => "001001111100001010111",
		320 => "001001111100001010111",
		321 => "001000000100101110110",
		322 => "001000000100101110110",
		323 => "001000000100101110110",
		324 => "011000000101111110011",
		325 => "011000000101111110011",
		326 => "011000000101111110011",
		327 => "011000101100111010001",
		328 => "011000101100111010001",
		329 => "011000101100111010001",
		330 => "001001111100001010111",
		331 => "001001111100001010111",
		332 => "001001111100001010111",
		333 => "001000000100101110110",
		334 => "001000000100101110110",
		335 => "001000000100101110110",
		336 => "011000000101111110011",
		337 => "011000000101111110011",
		338 => "011000000101111110011",
		339 => "011000101100111010001",
		340 => "011000101100111010001",
		341 => "011000101100111010001",
		342 => "001001111100001010111",
		343 => "001001111100001010111",
		344 => "001001111100001010111",
		345 => "001000000100101110110",
		346 => "001000000100101110110",
		347 => "001000000100101110110",
		348 => "011000000101111110011",
		349 => "011000000101111110011",
		350 => "011000000101111110011",
		351 => "011000101100111010001",
		352 => "011000101100111010001",
		353 => "011000101100111010001",
		354 => "001001111100001010111",
		355 => "001001111100001010111",
		356 => "001001111100001010111",
		357 => "001000000100101110110",
		358 => "001000000100101110110",
		359 => "001000000100101110110",
		360 => "011000000101111110011",
		361 => "011000000101111110011",
		362 => "011000000101111110011",
		363 => "011000101100111010001",
		364 => "011000101100111010001",
		365 => "011000101100111010001",
		366 => "001001111100001010111",
		367 => "001001111100001010111",
		368 => "001001111100001010111",
		369 => "001000000100101110110",
		370 => "001000000100101110110",
		371 => "001000000100101110110",
		372 => "011000000101111110011",
		373 => "011000000101111110011",
		374 => "011000000101111110011",
		375 => "011000101100111010001",
		376 => "011000101100111010001",
		377 => "011000101100111010001",
		378 => "001001111100001010111",
		379 => "001001111100001010111",
		380 => "001001111100001010111",
		381 => "001000000100101110110",
		382 => "001000000100101110110",
		383 => "001000000100101110110",
		384 => "011010100100001110100",
		385 => "011010100100001110100",
		386 => "011010100100001110100",
		387 => "011010100100001110100",
		388 => "011010100100001110100",
		389 => "011010100100001110100",
		390 => "011010100100001110100",
		391 => "011010100100001110100",
		392 => "011010100100001110100",
		393 => "011010100100001110100",
		394 => "011010100100001110100",
		395 => "011010100100001110100",
		396 => "011010100100001110100",
		397 => "011010100100001110100",
		398 => "011010100100001110100",
		399 => "011010100100001110100",
		400 => "011010100100001110100",
		401 => "011010100100001110100",
		402 => "011010100100001110100",
		403 => "011010100100001110100",
		404 => "011010100100001110100",
		405 => "011010100100001110100",
		406 => "011010100100001110100",
		407 => "011010100100001110100",
		408 => "011010100100001110100",
		409 => "011010100100001110100",
		410 => "011010100100001110100",
		411 => "011010100100001110100",
		412 => "011010100100001110100",
		413 => "011010100100001110100",
		414 => "011010100100001110100",
		415 => "011010100100001110100",
		416 => "011010100100001110100",
		417 => "011010100100001110100",
		418 => "011010100100001110100",
		419 => "011010100100001110100",
		420 => "011010100100001110100",
		421 => "011010100100001110100",
		422 => "011010100100001110100",
		423 => "011010100100001110100",
		424 => "011010100100001110100",
		425 => "011010100100001110100",
		426 => "011010100100001110100",
		427 => "011010100100001110100",
		428 => "011010100100001110100",
		429 => "011010100100001110100",
		430 => "011010100100001110100",
		431 => "011010100100001110100",
		432 => "011010100100001110100",
		433 => "011010100100001110100",
		434 => "011010100100001110100",
		435 => "011010100100001110100",
		436 => "011010100100001110100",
		437 => "011010100100001110100",
		438 => "011010100100001110100",
		439 => "011010100100001110100",
		440 => "011010100100001110100",
		441 => "011010100100001110100",
		442 => "011010100100001110100",
		443 => "011010100100001110100",
		444 => "011010100100001110100",
		445 => "011010100100001110100",
		446 => "011010100100001110100",
		447 => "011010100100001110100",
		448 => "011010100100001110100",
		449 => "011010100100001110100",
		450 => "011010100100001110100",
		451 => "011010100100001110100",
		452 => "011010100100001110100",
		453 => "011010100100001110100",
		454 => "011010100100001110100",
		455 => "011010100100001110100",
		456 => "011010100100001110100",
		457 => "011010100100001110100",
		458 => "011010100100001110100",
		459 => "011010100100001110100",
		460 => "011010100100001110100",
		461 => "011010100100001110100",
		462 => "011010100100001110100",
		463 => "011010100100001110100",
		464 => "011010100100001110100",
		465 => "011010100100001110100",
		466 => "011010100100001110100",
		467 => "011010100100001110100",
		468 => "011010100100001110100",
		469 => "011010100100001110100",
		470 => "011010100100001110100",
		471 => "011010100100001110100",
		472 => "011010100100001110100",
		473 => "011010100100001110100",
		474 => "011010100100001110100",
		475 => "011010100100001110100",
		476 => "011010100100001110100",
		477 => "011010100100001110100",
		478 => "011010100100001110100",
		479 => "011010100100001110100",
		480 => "011001111100001010110",
		481 => "011001111100001010110",
		482 => "011001111100001010110",
		483 => "011001111100001010110",
		484 => "011001111100001010110",
		485 => "011001111100001010110",
		486 => "011001111100001010110",
		487 => "011001111100001010110",
		488 => "011001111100001010110",
		489 => "011001111100001010110",
		490 => "011001111100001010110",
		491 => "011001111100001010110",
		492 => "011001111100001010110",
		493 => "011001111100001010110",
		494 => "011001111100001010110",
		495 => "011001111100001010110",
		496 => "011001111100001010110",
		497 => "011001111100001010110",
		498 => "011001111100001010110",
		499 => "011001111100001010110",
		500 => "011001111100001010110",
		501 => "011001111100001010110",
		502 => "011001111100001010110",
		503 => "011001111100001010110",
		504 => "011001111100001010110",
		505 => "011001111100001010110",
		506 => "011001111100001010110",
		507 => "011001111100001010110",
		508 => "011001111100001010110",
		509 => "011001111100001010110",
		510 => "011001111100001010110",
		511 => "011001111100001010110",
		512 => "011001111100001010110",
		513 => "011001111100001010110",
		514 => "011001111100001010110",
		515 => "011001111100001010110",
		516 => "011001111100001010110",
		517 => "011001111100001010110",
		518 => "011001111100001010110",
		519 => "011001111100001010110",
		520 => "011001111100001010110",
		521 => "011001111100001010110",
		522 => "011001111100001010110",
		523 => "011001111100001010110",
		524 => "011001111100001010110",
		525 => "011001111100001010110",
		526 => "011001111100001010110",
		527 => "011001111100001010110",
		528 => "011001111100001010110",
		529 => "011001111100001010110",
		530 => "011001111100001010110",
		531 => "011001111100001010110",
		532 => "011001111100001010110",
		533 => "011001111100001010110",
		534 => "011001111100001010110",
		535 => "011001111100001010110",
		536 => "011001111100001010110",
		537 => "011001111100001010110",
		538 => "011001111100001010110",
		539 => "011001111100001010110",
		540 => "011001111100001010110",
		541 => "011001111100001010110",
		542 => "011001111100001010110",
		543 => "011001111100001010110",
		544 => "011001111100001010110",
		545 => "011001111100001010110",
		546 => "011001111100001010110",
		547 => "011001111100001010110",
		548 => "011001111100001010110",
		549 => "011001111100001010110",
		550 => "011001111100001010110",
		551 => "011001111100001010110",
		552 => "011001111100001010110",
		553 => "011001111100001010110",
		554 => "011001111100001010110",
		555 => "011001111100001010110",
		556 => "011001111100001010110",
		557 => "011001111100001010110",
		558 => "011001111100001010110",
		559 => "011001111100001010110",
		560 => "011001111100001010110",
		561 => "011001111100001010110",
		562 => "011001111100001010110",
		563 => "011001111100001010110",
		564 => "011001111100001010110",
		565 => "011001111100001010110",
		566 => "011001111100001010110",
		567 => "011001111100001010110",
		568 => "011001111100001010110",
		569 => "011001111100001010110",
		570 => "011001111100001010110",
		571 => "011001111100001010110",
		572 => "011001111100001010110",
		573 => "011001111100001010110",
		574 => "011001111100001010110",
		575 => "011001111100001010110",
		576 => "011000101100100010101",
		577 => "011000101100100010101",
		578 => "011000101100100010101",
		579 => "011000101100100010101",
		580 => "011000101100100010101",
		581 => "011000101100100010101",
		582 => "011000101100100010101",
		583 => "011000101100100010101",
		584 => "011000101100100010101",
		585 => "011000101100100010101",
		586 => "011000101100100010101",
		587 => "011000101100100010101",
		588 => "011000101100100010101",
		589 => "011000101100100010101",
		590 => "011000101100100010101",
		591 => "011000101100100010101",
		592 => "011000101100100010101",
		593 => "011000101100100010101",
		594 => "011000101100100010101",
		595 => "011000101100100010101",
		596 => "011000101100100010101",
		597 => "011000101100100010101",
		598 => "011000101100100010101",
		599 => "011000101100100010101",
		600 => "011000101100100010101",
		601 => "011000101100100010101",
		602 => "011000101100100010101",
		603 => "011000101100100010101",
		604 => "011000101100100010101",
		605 => "011000101100100010101",
		606 => "011000101100100010101",
		607 => "011000101100100010101",
		608 => "011000101100100010101",
		609 => "011000101100100010101",
		610 => "011000101100100010101",
		611 => "011000101100100010101",
		612 => "011000101100100010101",
		613 => "011000101100100010101",
		614 => "011000101100100010101",
		615 => "011000101100100010101",
		616 => "011000101100100010101",
		617 => "011000101100100010101",
		618 => "011000101100100010101",
		619 => "011000101100100010101",
		620 => "011000101100100010101",
		621 => "011000101100100010101",
		622 => "011000101100100010101",
		623 => "011000101100100010101",
		624 => "011000101100100010101",
		625 => "011000101100100010101",
		626 => "011000101100100010101",
		627 => "011000101100100010101",
		628 => "011000101100100010101",
		629 => "011000101100100010101",
		630 => "011000101100100010101",
		631 => "011000101100100010101",
		632 => "011000101100100010101",
		633 => "011000101100100010101",
		634 => "011000101100100010101",
		635 => "011000101100100010101",
		636 => "011000101100100010101",
		637 => "011000101100100010101",
		638 => "011000101100100010101",
		639 => "011000101100100010101",
		640 => "011000101100100010101",
		641 => "011000101100100010101",
		642 => "011000101100100010101",
		643 => "011000101100100010101",
		644 => "011000101100100010101",
		645 => "011000101100100010101",
		646 => "011000101100100010101",
		647 => "011000101100100010101",
		648 => "011000101100100010101",
		649 => "011000101100100010101",
		650 => "011000101100100010101",
		651 => "011000101100100010101",
		652 => "011000101100100010101",
		653 => "011000101100100010101",
		654 => "011000101100100010101",
		655 => "011000101100100010101",
		656 => "011000101100100010101",
		657 => "011000101100100010101",
		658 => "011000101100100010101",
		659 => "011000101100100010101",
		660 => "011000101100100010101",
		661 => "011000101100100010101",
		662 => "011000101100100010101",
		663 => "011000101100100010101",
		664 => "011000101100100010101",
		665 => "011000101100100010101",
		666 => "011000101100100010101",
		667 => "011000101100100010101",
		668 => "011000101100100010101",
		669 => "011000101100100010101",
		670 => "011000101100100010101",
		671 => "011000101100100010101",
		672 => "011000101100100110010",
		673 => "011000101100100110010",
		674 => "011000101100100110010",
		675 => "011000101100100110010",
		676 => "011000101100100110010",
		677 => "011000101100100110010",
		678 => "011000101100100110010",
		679 => "011000101100100110010",
		680 => "011000101100100110010",
		681 => "011000101100100110010",
		682 => "011000101100100110010",
		683 => "011000101100100110010",
		684 => "011000101100100110010",
		685 => "011000101100100110010",
		686 => "011000101100100110010",
		687 => "011000101100100110010",
		688 => "011000101100100110010",
		689 => "011000101100100110010",
		690 => "011000101100100110010",
		691 => "011000101100100110010",
		692 => "011000101100100110010",
		693 => "011000101100100110010",
		694 => "011000101100100110010",
		695 => "011000101100100110010",
		696 => "011000101100100110010",
		697 => "011000101100100110010",
		698 => "011000101100100110010",
		699 => "011000101100100110010",
		700 => "011000101100100110010",
		701 => "011000101100100110010",
		702 => "011000101100100110010",
		703 => "011000101100100110010",
		704 => "011000101100100110010",
		705 => "011000101100100110010",
		706 => "011000101100100110010",
		707 => "011000101100100110010",
		708 => "011000101100100110010",
		709 => "011000101100100110010",
		710 => "011000101100100110010",
		711 => "011000101100100110010",
		712 => "011000101100100110010",
		713 => "011000101100100110010",
		714 => "011000101100100110010",
		715 => "011000101100100110010",
		716 => "011000101100100110010",
		717 => "011000101100100110010",
		718 => "011000101100100110010",
		719 => "011000101100100110010",
		720 => "011000101100100110010",
		721 => "011000101100100110010",
		722 => "011000101100100110010",
		723 => "011000101100100110010",
		724 => "011000101100100110010",
		725 => "011000101100100110010",
		726 => "011000101100100110010",
		727 => "011000101100100110010",
		728 => "011000101100100110010",
		729 => "011000101100100110010",
		730 => "011000101100100110010",
		731 => "011000101100100110010",
		732 => "011000101100100110010",
		733 => "011000101100100110010",
		734 => "011000101100100110010",
		735 => "011000101100100110010",
		736 => "011000101100100110010",
		737 => "011000101100100110010",
		738 => "011000101100100110010",
		739 => "011000101100100110010",
		740 => "011000101100100110010",
		741 => "011000101100100110010",
		742 => "011000101100100110010",
		743 => "011000101100100110010",
		744 => "011000101100100110010",
		745 => "011000101100100110010",
		746 => "011000101100100110010",
		747 => "011000101100100110010",
		748 => "011000101100100110010",
		749 => "011000101100100110010",
		750 => "011000101100100110010",
		751 => "011000101100100110010",
		752 => "011000101100100110010",
		753 => "011000101100100110010",
		754 => "011000101100100110010",
		755 => "011000101100100110010",
		756 => "011000101100100110010",
		757 => "011000101100100110010",
		758 => "011000101100100110010",
		759 => "011000101100100110010",
		760 => "011000101100100110010",
		761 => "011000101100100110010",
		762 => "011000101100100110010",
		763 => "011000101100100110010",
		764 => "011000101100100110010",
		765 => "011000101100100110010",
		766 => "011000101100100110010",
		767 => "011000101100100110010",
		768 => "111000010100001010000",
		769 => "111000010100001010000",
		770 => "111000010100001010000",
		771 => "111000010100001010000",
		772 => "111000010100001010000",
		773 => "111000010100001010000",
		774 => "111000010100001010000",
		775 => "111000010100001010000",
		776 => "111000010100001010000",
		777 => "111000010100001010000",
		778 => "111000010100001010000",
		779 => "111000010100001010000",
		780 => "111000010100001010000",
		781 => "111000010100001010000",
		782 => "111000010100001010000",
		783 => "111000010100001010000",
		784 => "111000010100001010000",
		785 => "111000010100001010000",
		786 => "111000010100001010000",
		787 => "111000010100001010000",
		788 => "111000010100001010000",
		789 => "111000010100001010000",
		790 => "111000010100001010000",
		791 => "111000010100001010000",
		792 => "111000010100001010000",
		793 => "111000010100001010000",
		794 => "111000010100001010000",
		795 => "111000010100001010000",
		796 => "111000010100001010000",
		797 => "111000010100001010000",
		798 => "111000010100001010000",
		799 => "111000010100001010000",
		800 => "111000010100001010000",
		801 => "111000010100001010000",
		802 => "111000010100001010000",
		803 => "111000010100001010000",
		804 => "111000010100001010000",
		805 => "111000010100001010000",
		806 => "111000010100001010000",
		807 => "111000010100001010000",
		808 => "111000010100001010000",
		809 => "111000010100001010000",
		810 => "111000010100001010000",
		811 => "111000010100001010000",
		812 => "111000010100001010000",
		813 => "111000010100001010000",
		814 => "111000010100001010000",
		815 => "111000010100001010000",
		816 => "111000010100001010000",
		817 => "111000010100001010000",
		818 => "111000010100001010000",
		819 => "111000010100001010000",
		820 => "111000010100001010000",
		821 => "111000010100001010000",
		822 => "111000010100001010000",
		823 => "111000010100001010000",
		824 => "111000010100001010000",
		825 => "111000010100001010000",
		826 => "111000010100001010000",
		827 => "111000010100001010000",
		828 => "111000010100001010000",
		829 => "111000010100001010000",
		830 => "111000010100001010000",
		831 => "111000010100001010000",
		832 => "111000010100001010000",
		833 => "111000010100001010000",
		834 => "111000010100001010000",
		835 => "111000010100001010000",
		836 => "111000010100001010000",
		837 => "111000010100001010000",
		838 => "111000010100001010000",
		839 => "111000010100001010000",
		840 => "111000010100001010000",
		841 => "111000010100001010000",
		842 => "111000010100001010000",
		843 => "111000010100001010000",
		844 => "111000010100001010000",
		845 => "111000010100001010000",
		846 => "111000010100001010000",
		847 => "111000010100001010000",
		848 => "111000010100001010000",
		849 => "111000010100001010000",
		850 => "111000010100001010000",
		851 => "111000010100001010000",
		852 => "111000010100001010000",
		853 => "111000010100001010000",
		854 => "111000010100001010000",
		855 => "111000010100001010000",
		856 => "111000010100001010000",
		857 => "111000010100001010000",
		858 => "111000010100001010000",
		859 => "111000010100001010000",
		860 => "111000010100001010000",
		861 => "111000010100001010000",
		862 => "111000010100001010000",
		863 => "111000010100001010000");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;