----------------------------------------------------------------------------------
--                                    The Mux
--
--   Sequential component for select each InputButterflySelectOut of butterfly.
--   
--   InputButterflySelectOut -- 
--   OutputButterfly -- 
--   Control -- Select InputButterfly
--
----------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_unsigned.ALL;
USE IEEE.numeric_std.ALL;
USE work.MainPackage.all;

ENTITY SelectOut IS
    GENERIC(NFFT : INTEGER);
    PORT(
        ControlSelectOut : IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
        InputSelectOut : IN ComplexVector((NFFT-1) DOWNTO 0);
        OutputSelectOut : OUT ComplexVector((NFFT-1) DOWNTO 0)
        );
END SelectOut;

ARCHITECTURE Behavioral OF SelectOut IS

BEGIN

OutputSelectOut(0) <= InputSelectOut(0);
OutputSelectOut(1) <= InputSelectOut(256) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(256) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(128) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(64) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(32) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(16) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(8) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(4) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(2);
OutputSelectOut(2) <= InputSelectOut(1) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(2) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(2) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(2) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(2) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(2) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(2) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(2) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(1);
OutputSelectOut(3) <= InputSelectOut(257) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(258) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(130) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(66) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(34) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(18) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(10) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(6) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(3);
OutputSelectOut(4) <= InputSelectOut(2) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(4) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(4) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(4) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(4) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(4) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(4) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(1) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(4);
OutputSelectOut(5) <= InputSelectOut(258) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(260) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(132) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(68) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(36) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(20) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(12) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(5) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(6);
OutputSelectOut(6) <= InputSelectOut(3) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(6) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(6) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(6) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(6) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(6) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(6) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(3) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(5);
OutputSelectOut(7) <= InputSelectOut(259) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(262) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(134) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(70) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(38) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(22) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(14) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(7) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(7);
OutputSelectOut(8) <= InputSelectOut(4) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(8) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(8) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(8) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(8) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(8) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(1) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(8) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(8);
OutputSelectOut(9) <= InputSelectOut(260) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(264) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(136) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(72) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(40) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(24) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(9) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(12) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(10);
OutputSelectOut(10) <= InputSelectOut(5) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(10) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(10) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(10) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(10) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(10) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(3) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(10) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(9);
OutputSelectOut(11) <= InputSelectOut(261) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(266) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(138) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(74) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(42) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(26) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(11) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(14) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(11);
OutputSelectOut(12) <= InputSelectOut(6) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(12) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(12) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(12) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(12) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(12) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(5) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(9) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(12);
OutputSelectOut(13) <= InputSelectOut(262) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(268) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(140) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(76) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(44) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(28) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(13) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(13) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(14);
OutputSelectOut(14) <= InputSelectOut(7) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(14) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(14) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(14) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(14) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(14) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(7) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(11) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(13);
OutputSelectOut(15) <= InputSelectOut(263) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(270) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(142) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(78) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(46) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(30) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(15) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(15) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(15);
OutputSelectOut(16) <= InputSelectOut(8) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(16) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(16) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(16) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(16) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(1) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(16) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(16) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(16);
OutputSelectOut(17) <= InputSelectOut(264) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(272) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(144) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(80) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(48) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(17) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(24) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(20) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(18);
OutputSelectOut(18) <= InputSelectOut(9) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(18) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(18) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(18) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(18) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(3) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(18) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(18) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(17);
OutputSelectOut(19) <= InputSelectOut(265) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(274) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(146) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(82) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(50) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(19) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(26) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(22) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(19);
OutputSelectOut(20) <= InputSelectOut(10) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(20) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(20) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(20) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(20) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(5) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(20) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(17) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(20);
OutputSelectOut(21) <= InputSelectOut(266) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(276) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(148) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(84) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(52) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(21) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(28) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(21) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(22);
OutputSelectOut(22) <= InputSelectOut(11) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(22) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(22) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(22) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(22) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(7) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(22) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(19) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(21);
OutputSelectOut(23) <= InputSelectOut(267) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(278) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(150) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(86) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(54) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(23) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(30) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(23) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(23);
OutputSelectOut(24) <= InputSelectOut(12) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(24) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(24) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(24) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(24) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(9) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(17) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(24) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(24);
OutputSelectOut(25) <= InputSelectOut(268) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(280) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(152) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(88) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(56) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(25) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(25) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(28) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(26);
OutputSelectOut(26) <= InputSelectOut(13) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(26) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(26) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(26) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(26) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(11) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(19) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(26) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(25);
OutputSelectOut(27) <= InputSelectOut(269) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(282) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(154) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(90) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(58) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(27) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(27) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(30) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(27);
OutputSelectOut(28) <= InputSelectOut(14) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(28) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(28) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(28) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(28) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(13) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(21) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(25) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(28);
OutputSelectOut(29) <= InputSelectOut(270) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(284) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(156) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(92) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(60) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(29) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(29) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(29) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(30);
OutputSelectOut(30) <= InputSelectOut(15) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(30) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(30) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(30) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(30) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(15) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(23) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(27) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(29);
OutputSelectOut(31) <= InputSelectOut(271) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(286) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(158) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(94) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(62) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(31) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(31) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(31) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(31);
OutputSelectOut(32) <= InputSelectOut(16) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(32) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(32) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(32) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(1) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(32) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(32) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(32) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(32);
OutputSelectOut(33) <= InputSelectOut(272) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(288) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(160) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(96) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(33) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(48) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(40) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(36) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(34);
OutputSelectOut(34) <= InputSelectOut(17) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(34) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(34) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(34) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(3) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(34) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(34) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(34) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(33);
OutputSelectOut(35) <= InputSelectOut(273) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(290) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(162) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(98) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(35) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(50) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(42) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(38) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(35);
OutputSelectOut(36) <= InputSelectOut(18) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(36) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(36) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(36) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(5) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(36) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(36) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(33) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(36);
OutputSelectOut(37) <= InputSelectOut(274) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(292) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(164) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(100) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(37) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(52) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(44) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(37) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(38);
OutputSelectOut(38) <= InputSelectOut(19) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(38) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(38) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(38) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(7) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(38) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(38) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(35) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(37);
OutputSelectOut(39) <= InputSelectOut(275) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(294) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(166) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(102) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(39) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(54) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(46) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(39) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(39);
OutputSelectOut(40) <= InputSelectOut(20) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(40) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(40) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(40) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(9) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(40) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(33) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(40) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(40);
OutputSelectOut(41) <= InputSelectOut(276) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(296) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(168) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(104) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(41) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(56) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(41) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(44) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(42);
OutputSelectOut(42) <= InputSelectOut(21) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(42) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(42) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(42) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(11) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(42) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(35) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(42) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(41);
OutputSelectOut(43) <= InputSelectOut(277) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(298) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(170) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(106) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(43) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(58) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(43) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(46) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(43);
OutputSelectOut(44) <= InputSelectOut(22) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(44) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(44) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(44) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(13) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(44) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(37) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(41) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(44);
OutputSelectOut(45) <= InputSelectOut(278) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(300) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(172) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(108) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(45) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(60) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(45) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(45) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(46);
OutputSelectOut(46) <= InputSelectOut(23) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(46) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(46) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(46) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(15) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(46) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(39) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(43) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(45);
OutputSelectOut(47) <= InputSelectOut(279) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(302) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(174) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(110) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(47) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(62) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(47) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(47) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(47);
OutputSelectOut(48) <= InputSelectOut(24) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(48) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(48) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(48) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(17) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(33) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(48) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(48) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(48);
OutputSelectOut(49) <= InputSelectOut(280) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(304) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(176) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(112) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(49) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(49) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(56) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(52) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(50);
OutputSelectOut(50) <= InputSelectOut(25) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(50) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(50) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(50) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(19) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(35) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(50) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(50) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(49);
OutputSelectOut(51) <= InputSelectOut(281) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(306) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(178) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(114) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(51) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(51) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(58) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(54) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(51);
OutputSelectOut(52) <= InputSelectOut(26) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(52) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(52) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(52) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(21) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(37) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(52) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(49) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(52);
OutputSelectOut(53) <= InputSelectOut(282) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(308) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(180) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(116) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(53) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(53) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(60) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(53) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(54);
OutputSelectOut(54) <= InputSelectOut(27) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(54) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(54) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(54) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(23) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(39) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(54) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(51) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(53);
OutputSelectOut(55) <= InputSelectOut(283) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(310) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(182) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(118) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(55) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(55) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(62) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(55) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(55);
OutputSelectOut(56) <= InputSelectOut(28) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(56) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(56) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(56) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(25) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(41) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(49) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(56) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(56);
OutputSelectOut(57) <= InputSelectOut(284) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(312) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(184) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(120) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(57) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(57) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(57) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(60) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(58);
OutputSelectOut(58) <= InputSelectOut(29) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(58) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(58) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(58) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(27) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(43) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(51) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(58) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(57);
OutputSelectOut(59) <= InputSelectOut(285) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(314) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(186) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(122) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(59) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(59) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(59) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(62) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(59);
OutputSelectOut(60) <= InputSelectOut(30) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(60) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(60) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(60) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(29) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(45) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(53) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(57) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(60);
OutputSelectOut(61) <= InputSelectOut(286) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(316) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(188) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(124) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(61) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(61) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(61) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(61) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(62);
OutputSelectOut(62) <= InputSelectOut(31) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(62) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(62) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(62) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(31) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(47) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(55) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(59) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(61);
OutputSelectOut(63) <= InputSelectOut(287) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(318) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(190) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(126) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(63) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(63) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(63) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(63) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(63);
OutputSelectOut(64) <= InputSelectOut(32) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(64) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(64) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(1) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(64) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(64) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(64) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(64) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(64);
OutputSelectOut(65) <= InputSelectOut(288) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(320) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(192) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(65) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(96) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(80) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(72) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(68) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(66);
OutputSelectOut(66) <= InputSelectOut(33) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(66) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(66) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(3) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(66) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(66) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(66) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(66) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(65);
OutputSelectOut(67) <= InputSelectOut(289) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(322) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(194) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(67) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(98) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(82) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(74) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(70) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(67);
OutputSelectOut(68) <= InputSelectOut(34) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(68) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(68) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(5) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(68) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(68) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(68) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(65) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(68);
OutputSelectOut(69) <= InputSelectOut(290) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(324) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(196) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(69) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(100) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(84) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(76) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(69) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(70);
OutputSelectOut(70) <= InputSelectOut(35) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(70) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(70) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(7) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(70) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(70) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(70) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(67) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(69);
OutputSelectOut(71) <= InputSelectOut(291) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(326) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(198) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(71) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(102) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(86) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(78) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(71) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(71);
OutputSelectOut(72) <= InputSelectOut(36) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(72) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(72) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(9) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(72) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(72) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(65) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(72) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(72);
OutputSelectOut(73) <= InputSelectOut(292) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(328) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(200) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(73) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(104) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(88) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(73) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(76) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(74);
OutputSelectOut(74) <= InputSelectOut(37) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(74) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(74) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(11) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(74) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(74) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(67) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(74) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(73);
OutputSelectOut(75) <= InputSelectOut(293) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(330) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(202) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(75) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(106) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(90) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(75) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(78) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(75);
OutputSelectOut(76) <= InputSelectOut(38) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(76) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(76) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(13) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(76) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(76) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(69) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(73) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(76);
OutputSelectOut(77) <= InputSelectOut(294) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(332) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(204) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(77) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(108) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(92) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(77) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(77) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(78);
OutputSelectOut(78) <= InputSelectOut(39) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(78) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(78) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(15) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(78) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(78) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(71) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(75) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(77);
OutputSelectOut(79) <= InputSelectOut(295) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(334) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(206) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(79) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(110) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(94) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(79) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(79) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(79);
OutputSelectOut(80) <= InputSelectOut(40) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(80) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(80) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(17) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(80) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(65) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(80) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(80) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(80);
OutputSelectOut(81) <= InputSelectOut(296) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(336) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(208) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(81) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(112) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(81) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(88) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(84) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(82);
OutputSelectOut(82) <= InputSelectOut(41) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(82) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(82) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(19) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(82) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(67) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(82) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(82) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(81);
OutputSelectOut(83) <= InputSelectOut(297) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(338) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(210) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(83) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(114) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(83) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(90) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(86) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(83);
OutputSelectOut(84) <= InputSelectOut(42) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(84) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(84) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(21) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(84) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(69) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(84) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(81) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(84);
OutputSelectOut(85) <= InputSelectOut(298) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(340) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(212) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(85) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(116) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(85) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(92) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(85) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(86);
OutputSelectOut(86) <= InputSelectOut(43) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(86) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(86) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(23) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(86) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(71) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(86) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(83) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(85);
OutputSelectOut(87) <= InputSelectOut(299) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(342) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(214) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(87) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(118) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(87) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(94) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(87) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(87);
OutputSelectOut(88) <= InputSelectOut(44) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(88) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(88) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(25) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(88) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(73) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(81) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(88) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(88);
OutputSelectOut(89) <= InputSelectOut(300) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(344) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(216) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(89) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(120) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(89) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(89) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(92) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(90);
OutputSelectOut(90) <= InputSelectOut(45) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(90) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(90) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(27) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(90) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(75) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(83) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(90) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(89);
OutputSelectOut(91) <= InputSelectOut(301) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(346) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(218) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(91) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(122) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(91) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(91) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(94) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(91);
OutputSelectOut(92) <= InputSelectOut(46) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(92) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(92) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(29) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(92) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(77) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(85) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(89) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(92);
OutputSelectOut(93) <= InputSelectOut(302) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(348) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(220) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(93) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(124) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(93) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(93) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(93) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(94);
OutputSelectOut(94) <= InputSelectOut(47) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(94) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(94) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(31) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(94) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(79) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(87) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(91) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(93);
OutputSelectOut(95) <= InputSelectOut(303) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(350) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(222) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(95) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(126) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(95) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(95) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(95) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(95);
OutputSelectOut(96) <= InputSelectOut(48) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(96) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(96) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(33) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(65) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(96) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(96) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(96) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(96);
OutputSelectOut(97) <= InputSelectOut(304) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(352) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(224) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(97) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(97) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(112) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(104) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(100) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(98);
OutputSelectOut(98) <= InputSelectOut(49) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(98) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(98) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(35) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(67) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(98) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(98) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(98) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(97);
OutputSelectOut(99) <= InputSelectOut(305) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(354) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(226) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(99) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(99) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(114) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(106) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(102) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(99);
OutputSelectOut(100) <= InputSelectOut(50) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(100) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(100) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(37) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(69) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(100) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(100) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(97) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(100);
OutputSelectOut(101) <= InputSelectOut(306) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(356) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(228) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(101) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(101) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(116) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(108) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(101) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(102);
OutputSelectOut(102) <= InputSelectOut(51) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(102) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(102) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(39) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(71) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(102) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(102) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(99) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(101);
OutputSelectOut(103) <= InputSelectOut(307) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(358) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(230) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(103) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(103) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(118) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(110) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(103) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(103);
OutputSelectOut(104) <= InputSelectOut(52) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(104) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(104) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(41) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(73) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(104) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(97) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(104) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(104);
OutputSelectOut(105) <= InputSelectOut(308) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(360) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(232) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(105) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(105) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(120) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(105) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(108) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(106);
OutputSelectOut(106) <= InputSelectOut(53) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(106) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(106) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(43) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(75) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(106) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(99) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(106) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(105);
OutputSelectOut(107) <= InputSelectOut(309) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(362) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(234) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(107) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(107) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(122) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(107) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(110) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(107);
OutputSelectOut(108) <= InputSelectOut(54) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(108) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(108) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(45) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(77) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(108) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(101) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(105) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(108);
OutputSelectOut(109) <= InputSelectOut(310) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(364) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(236) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(109) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(109) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(124) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(109) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(109) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(110);
OutputSelectOut(110) <= InputSelectOut(55) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(110) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(110) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(47) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(79) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(110) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(103) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(107) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(109);
OutputSelectOut(111) <= InputSelectOut(311) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(366) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(238) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(111) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(111) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(126) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(111) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(111) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(111);
OutputSelectOut(112) <= InputSelectOut(56) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(112) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(112) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(49) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(81) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(97) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(112) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(112) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(112);
OutputSelectOut(113) <= InputSelectOut(312) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(368) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(240) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(113) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(113) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(113) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(120) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(116) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(114);
OutputSelectOut(114) <= InputSelectOut(57) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(114) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(114) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(51) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(83) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(99) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(114) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(114) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(113);
OutputSelectOut(115) <= InputSelectOut(313) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(370) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(242) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(115) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(115) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(115) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(122) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(118) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(115);
OutputSelectOut(116) <= InputSelectOut(58) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(116) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(116) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(53) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(85) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(101) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(116) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(113) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(116);
OutputSelectOut(117) <= InputSelectOut(314) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(372) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(244) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(117) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(117) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(117) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(124) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(117) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(118);
OutputSelectOut(118) <= InputSelectOut(59) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(118) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(118) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(55) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(87) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(103) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(118) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(115) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(117);
OutputSelectOut(119) <= InputSelectOut(315) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(374) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(246) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(119) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(119) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(119) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(126) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(119) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(119);
OutputSelectOut(120) <= InputSelectOut(60) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(120) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(120) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(57) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(89) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(105) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(113) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(120) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(120);
OutputSelectOut(121) <= InputSelectOut(316) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(376) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(248) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(121) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(121) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(121) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(121) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(124) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(122);
OutputSelectOut(122) <= InputSelectOut(61) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(122) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(122) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(59) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(91) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(107) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(115) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(122) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(121);
OutputSelectOut(123) <= InputSelectOut(317) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(378) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(250) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(123) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(123) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(123) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(123) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(126) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(123);
OutputSelectOut(124) <= InputSelectOut(62) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(124) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(124) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(61) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(93) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(109) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(117) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(121) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(124);
OutputSelectOut(125) <= InputSelectOut(318) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(380) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(252) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(125) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(125) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(125) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(125) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(125) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(126);
OutputSelectOut(126) <= InputSelectOut(63) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(126) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(126) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(63) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(95) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(111) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(119) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(123) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(125);
OutputSelectOut(127) <= InputSelectOut(319) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(382) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(254) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(127) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(127) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(127) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(127) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(127) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(127);
OutputSelectOut(128) <= InputSelectOut(64) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(128) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(1) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(128) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(128) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(128) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(128) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(128) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(128);
OutputSelectOut(129) <= InputSelectOut(320) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(384) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(129) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(192) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(160) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(144) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(136) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(132) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(130);
OutputSelectOut(130) <= InputSelectOut(65) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(130) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(3) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(130) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(130) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(130) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(130) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(130) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(129);
OutputSelectOut(131) <= InputSelectOut(321) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(386) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(131) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(194) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(162) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(146) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(138) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(134) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(131);
OutputSelectOut(132) <= InputSelectOut(66) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(132) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(5) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(132) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(132) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(132) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(132) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(129) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(132);
OutputSelectOut(133) <= InputSelectOut(322) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(388) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(133) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(196) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(164) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(148) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(140) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(133) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(134);
OutputSelectOut(134) <= InputSelectOut(67) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(134) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(7) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(134) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(134) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(134) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(134) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(131) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(133);
OutputSelectOut(135) <= InputSelectOut(323) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(390) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(135) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(198) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(166) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(150) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(142) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(135) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(135);
OutputSelectOut(136) <= InputSelectOut(68) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(136) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(9) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(136) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(136) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(136) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(129) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(136) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(136);
OutputSelectOut(137) <= InputSelectOut(324) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(392) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(137) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(200) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(168) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(152) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(137) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(140) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(138);
OutputSelectOut(138) <= InputSelectOut(69) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(138) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(11) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(138) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(138) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(138) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(131) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(138) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(137);
OutputSelectOut(139) <= InputSelectOut(325) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(394) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(139) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(202) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(170) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(154) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(139) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(142) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(139);
OutputSelectOut(140) <= InputSelectOut(70) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(140) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(13) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(140) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(140) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(140) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(133) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(137) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(140);
OutputSelectOut(141) <= InputSelectOut(326) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(396) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(141) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(204) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(172) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(156) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(141) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(141) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(142);
OutputSelectOut(142) <= InputSelectOut(71) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(142) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(15) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(142) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(142) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(142) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(135) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(139) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(141);
OutputSelectOut(143) <= InputSelectOut(327) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(398) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(143) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(206) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(174) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(158) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(143) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(143) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(143);
OutputSelectOut(144) <= InputSelectOut(72) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(144) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(17) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(144) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(144) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(129) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(144) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(144) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(144);
OutputSelectOut(145) <= InputSelectOut(328) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(400) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(145) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(208) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(176) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(145) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(152) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(148) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(146);
OutputSelectOut(146) <= InputSelectOut(73) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(146) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(19) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(146) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(146) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(131) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(146) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(146) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(145);
OutputSelectOut(147) <= InputSelectOut(329) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(402) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(147) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(210) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(178) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(147) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(154) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(150) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(147);
OutputSelectOut(148) <= InputSelectOut(74) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(148) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(21) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(148) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(148) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(133) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(148) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(145) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(148);
OutputSelectOut(149) <= InputSelectOut(330) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(404) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(149) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(212) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(180) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(149) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(156) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(149) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(150);
OutputSelectOut(150) <= InputSelectOut(75) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(150) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(23) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(150) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(150) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(135) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(150) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(147) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(149);
OutputSelectOut(151) <= InputSelectOut(331) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(406) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(151) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(214) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(182) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(151) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(158) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(151) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(151);
OutputSelectOut(152) <= InputSelectOut(76) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(152) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(25) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(152) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(152) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(137) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(145) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(152) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(152);
OutputSelectOut(153) <= InputSelectOut(332) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(408) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(153) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(216) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(184) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(153) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(153) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(156) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(154);
OutputSelectOut(154) <= InputSelectOut(77) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(154) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(27) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(154) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(154) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(139) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(147) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(154) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(153);
OutputSelectOut(155) <= InputSelectOut(333) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(410) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(155) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(218) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(186) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(155) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(155) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(158) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(155);
OutputSelectOut(156) <= InputSelectOut(78) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(156) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(29) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(156) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(156) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(141) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(149) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(153) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(156);
OutputSelectOut(157) <= InputSelectOut(334) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(412) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(157) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(220) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(188) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(157) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(157) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(157) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(158);
OutputSelectOut(158) <= InputSelectOut(79) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(158) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(31) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(158) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(158) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(143) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(151) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(155) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(157);
OutputSelectOut(159) <= InputSelectOut(335) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(414) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(159) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(222) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(190) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(159) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(159) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(159) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(159);
OutputSelectOut(160) <= InputSelectOut(80) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(160) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(33) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(160) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(129) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(160) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(160) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(160) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(160);
OutputSelectOut(161) <= InputSelectOut(336) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(416) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(161) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(224) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(161) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(176) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(168) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(164) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(162);
OutputSelectOut(162) <= InputSelectOut(81) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(162) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(35) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(162) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(131) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(162) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(162) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(162) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(161);
OutputSelectOut(163) <= InputSelectOut(337) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(418) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(163) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(226) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(163) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(178) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(170) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(166) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(163);
OutputSelectOut(164) <= InputSelectOut(82) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(164) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(37) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(164) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(133) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(164) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(164) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(161) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(164);
OutputSelectOut(165) <= InputSelectOut(338) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(420) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(165) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(228) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(165) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(180) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(172) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(165) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(166);
OutputSelectOut(166) <= InputSelectOut(83) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(166) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(39) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(166) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(135) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(166) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(166) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(163) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(165);
OutputSelectOut(167) <= InputSelectOut(339) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(422) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(167) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(230) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(167) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(182) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(174) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(167) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(167);
OutputSelectOut(168) <= InputSelectOut(84) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(168) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(41) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(168) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(137) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(168) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(161) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(168) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(168);
OutputSelectOut(169) <= InputSelectOut(340) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(424) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(169) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(232) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(169) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(184) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(169) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(172) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(170);
OutputSelectOut(170) <= InputSelectOut(85) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(170) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(43) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(170) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(139) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(170) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(163) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(170) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(169);
OutputSelectOut(171) <= InputSelectOut(341) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(426) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(171) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(234) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(171) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(186) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(171) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(174) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(171);
OutputSelectOut(172) <= InputSelectOut(86) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(172) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(45) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(172) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(141) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(172) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(165) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(169) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(172);
OutputSelectOut(173) <= InputSelectOut(342) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(428) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(173) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(236) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(173) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(188) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(173) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(173) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(174);
OutputSelectOut(174) <= InputSelectOut(87) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(174) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(47) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(174) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(143) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(174) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(167) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(171) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(173);
OutputSelectOut(175) <= InputSelectOut(343) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(430) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(175) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(238) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(175) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(190) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(175) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(175) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(175);
OutputSelectOut(176) <= InputSelectOut(88) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(176) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(49) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(176) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(145) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(161) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(176) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(176) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(176);
OutputSelectOut(177) <= InputSelectOut(344) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(432) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(177) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(240) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(177) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(177) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(184) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(180) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(178);
OutputSelectOut(178) <= InputSelectOut(89) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(178) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(51) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(178) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(147) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(163) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(178) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(178) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(177);
OutputSelectOut(179) <= InputSelectOut(345) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(434) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(179) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(242) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(179) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(179) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(186) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(182) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(179);
OutputSelectOut(180) <= InputSelectOut(90) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(180) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(53) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(180) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(149) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(165) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(180) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(177) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(180);
OutputSelectOut(181) <= InputSelectOut(346) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(436) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(181) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(244) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(181) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(181) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(188) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(181) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(182);
OutputSelectOut(182) <= InputSelectOut(91) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(182) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(55) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(182) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(151) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(167) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(182) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(179) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(181);
OutputSelectOut(183) <= InputSelectOut(347) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(438) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(183) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(246) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(183) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(183) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(190) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(183) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(183);
OutputSelectOut(184) <= InputSelectOut(92) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(184) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(57) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(184) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(153) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(169) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(177) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(184) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(184);
OutputSelectOut(185) <= InputSelectOut(348) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(440) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(185) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(248) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(185) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(185) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(185) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(188) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(186);
OutputSelectOut(186) <= InputSelectOut(93) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(186) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(59) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(186) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(155) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(171) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(179) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(186) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(185);
OutputSelectOut(187) <= InputSelectOut(349) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(442) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(187) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(250) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(187) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(187) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(187) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(190) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(187);
OutputSelectOut(188) <= InputSelectOut(94) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(188) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(61) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(188) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(157) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(173) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(181) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(185) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(188);
OutputSelectOut(189) <= InputSelectOut(350) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(444) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(189) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(252) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(189) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(189) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(189) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(189) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(190);
OutputSelectOut(190) <= InputSelectOut(95) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(190) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(63) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(190) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(159) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(175) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(183) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(187) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(189);
OutputSelectOut(191) <= InputSelectOut(351) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(446) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(191) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(254) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(191) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(191) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(191) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(191) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(191);
OutputSelectOut(192) <= InputSelectOut(96) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(192) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(65) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(129) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(192) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(192) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(192) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(192) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(192);
OutputSelectOut(193) <= InputSelectOut(352) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(448) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(193) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(193) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(224) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(208) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(200) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(196) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(194);
OutputSelectOut(194) <= InputSelectOut(97) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(194) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(67) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(131) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(194) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(194) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(194) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(194) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(193);
OutputSelectOut(195) <= InputSelectOut(353) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(450) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(195) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(195) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(226) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(210) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(202) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(198) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(195);
OutputSelectOut(196) <= InputSelectOut(98) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(196) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(69) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(133) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(196) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(196) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(196) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(193) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(196);
OutputSelectOut(197) <= InputSelectOut(354) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(452) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(197) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(197) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(228) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(212) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(204) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(197) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(198);
OutputSelectOut(198) <= InputSelectOut(99) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(198) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(71) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(135) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(198) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(198) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(198) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(195) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(197);
OutputSelectOut(199) <= InputSelectOut(355) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(454) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(199) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(199) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(230) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(214) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(206) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(199) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(199);
OutputSelectOut(200) <= InputSelectOut(100) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(200) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(73) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(137) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(200) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(200) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(193) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(200) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(200);
OutputSelectOut(201) <= InputSelectOut(356) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(456) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(201) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(201) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(232) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(216) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(201) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(204) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(202);
OutputSelectOut(202) <= InputSelectOut(101) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(202) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(75) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(139) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(202) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(202) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(195) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(202) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(201);
OutputSelectOut(203) <= InputSelectOut(357) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(458) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(203) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(203) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(234) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(218) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(203) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(206) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(203);
OutputSelectOut(204) <= InputSelectOut(102) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(204) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(77) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(141) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(204) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(204) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(197) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(201) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(204);
OutputSelectOut(205) <= InputSelectOut(358) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(460) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(205) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(205) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(236) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(220) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(205) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(205) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(206);
OutputSelectOut(206) <= InputSelectOut(103) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(206) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(79) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(143) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(206) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(206) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(199) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(203) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(205);
OutputSelectOut(207) <= InputSelectOut(359) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(462) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(207) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(207) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(238) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(222) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(207) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(207) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(207);
OutputSelectOut(208) <= InputSelectOut(104) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(208) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(81) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(145) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(208) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(193) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(208) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(208) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(208);
OutputSelectOut(209) <= InputSelectOut(360) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(464) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(209) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(209) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(240) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(209) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(216) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(212) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(210);
OutputSelectOut(210) <= InputSelectOut(105) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(210) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(83) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(147) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(210) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(195) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(210) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(210) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(209);
OutputSelectOut(211) <= InputSelectOut(361) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(466) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(211) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(211) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(242) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(211) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(218) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(214) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(211);
OutputSelectOut(212) <= InputSelectOut(106) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(212) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(85) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(149) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(212) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(197) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(212) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(209) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(212);
OutputSelectOut(213) <= InputSelectOut(362) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(468) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(213) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(213) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(244) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(213) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(220) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(213) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(214);
OutputSelectOut(214) <= InputSelectOut(107) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(214) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(87) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(151) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(214) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(199) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(214) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(211) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(213);
OutputSelectOut(215) <= InputSelectOut(363) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(470) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(215) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(215) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(246) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(215) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(222) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(215) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(215);
OutputSelectOut(216) <= InputSelectOut(108) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(216) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(89) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(153) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(216) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(201) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(209) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(216) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(216);
OutputSelectOut(217) <= InputSelectOut(364) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(472) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(217) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(217) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(248) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(217) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(217) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(220) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(218);
OutputSelectOut(218) <= InputSelectOut(109) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(218) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(91) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(155) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(218) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(203) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(211) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(218) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(217);
OutputSelectOut(219) <= InputSelectOut(365) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(474) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(219) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(219) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(250) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(219) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(219) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(222) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(219);
OutputSelectOut(220) <= InputSelectOut(110) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(220) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(93) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(157) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(220) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(205) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(213) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(217) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(220);
OutputSelectOut(221) <= InputSelectOut(366) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(476) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(221) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(221) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(252) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(221) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(221) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(221) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(222);
OutputSelectOut(222) <= InputSelectOut(111) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(222) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(95) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(159) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(222) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(207) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(215) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(219) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(221);
OutputSelectOut(223) <= InputSelectOut(367) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(478) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(223) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(223) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(254) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(223) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(223) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(223) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(223);
OutputSelectOut(224) <= InputSelectOut(112) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(224) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(97) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(161) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(193) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(224) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(224) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(224) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(224);
OutputSelectOut(225) <= InputSelectOut(368) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(480) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(225) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(225) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(225) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(240) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(232) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(228) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(226);
OutputSelectOut(226) <= InputSelectOut(113) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(226) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(99) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(163) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(195) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(226) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(226) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(226) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(225);
OutputSelectOut(227) <= InputSelectOut(369) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(482) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(227) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(227) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(227) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(242) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(234) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(230) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(227);
OutputSelectOut(228) <= InputSelectOut(114) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(228) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(101) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(165) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(197) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(228) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(228) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(225) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(228);
OutputSelectOut(229) <= InputSelectOut(370) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(484) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(229) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(229) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(229) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(244) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(236) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(229) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(230);
OutputSelectOut(230) <= InputSelectOut(115) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(230) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(103) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(167) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(199) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(230) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(230) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(227) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(229);
OutputSelectOut(231) <= InputSelectOut(371) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(486) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(231) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(231) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(231) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(246) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(238) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(231) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(231);
OutputSelectOut(232) <= InputSelectOut(116) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(232) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(105) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(169) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(201) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(232) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(225) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(232) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(232);
OutputSelectOut(233) <= InputSelectOut(372) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(488) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(233) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(233) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(233) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(248) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(233) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(236) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(234);
OutputSelectOut(234) <= InputSelectOut(117) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(234) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(107) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(171) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(203) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(234) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(227) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(234) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(233);
OutputSelectOut(235) <= InputSelectOut(373) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(490) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(235) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(235) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(235) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(250) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(235) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(238) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(235);
OutputSelectOut(236) <= InputSelectOut(118) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(236) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(109) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(173) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(205) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(236) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(229) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(233) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(236);
OutputSelectOut(237) <= InputSelectOut(374) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(492) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(237) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(237) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(237) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(252) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(237) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(237) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(238);
OutputSelectOut(238) <= InputSelectOut(119) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(238) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(111) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(175) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(207) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(238) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(231) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(235) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(237);
OutputSelectOut(239) <= InputSelectOut(375) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(494) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(239) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(239) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(239) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(254) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(239) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(239) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(239);
OutputSelectOut(240) <= InputSelectOut(120) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(240) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(113) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(177) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(209) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(225) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(240) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(240) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(240);
OutputSelectOut(241) <= InputSelectOut(376) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(496) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(241) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(241) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(241) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(241) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(248) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(244) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(242);
OutputSelectOut(242) <= InputSelectOut(121) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(242) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(115) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(179) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(211) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(227) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(242) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(242) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(241);
OutputSelectOut(243) <= InputSelectOut(377) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(498) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(243) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(243) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(243) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(243) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(250) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(246) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(243);
OutputSelectOut(244) <= InputSelectOut(122) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(244) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(117) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(181) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(213) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(229) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(244) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(241) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(244);
OutputSelectOut(245) <= InputSelectOut(378) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(500) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(245) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(245) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(245) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(245) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(252) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(245) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(246);
OutputSelectOut(246) <= InputSelectOut(123) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(246) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(119) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(183) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(215) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(231) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(246) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(243) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(245);
OutputSelectOut(247) <= InputSelectOut(379) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(502) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(247) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(247) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(247) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(247) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(254) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(247) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(247);
OutputSelectOut(248) <= InputSelectOut(124) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(248) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(121) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(185) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(217) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(233) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(241) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(248) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(248);
OutputSelectOut(249) <= InputSelectOut(380) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(504) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(249) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(249) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(249) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(249) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(249) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(252) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(250);
OutputSelectOut(250) <= InputSelectOut(125) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(250) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(123) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(187) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(219) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(235) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(243) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(250) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(249);
OutputSelectOut(251) <= InputSelectOut(381) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(506) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(251) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(251) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(251) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(251) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(251) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(254) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(251);
OutputSelectOut(252) <= InputSelectOut(126) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(252) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(125) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(189) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(221) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(237) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(245) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(249) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(252);
OutputSelectOut(253) <= InputSelectOut(382) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(508) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(253) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(253) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(253) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(253) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(253) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(253) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(254);
OutputSelectOut(254) <= InputSelectOut(127) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(254) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(127) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(191) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(223) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(239) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(247) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(251) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(253);
OutputSelectOut(255) <= InputSelectOut(383) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(510) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(255) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(255) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(255) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(255) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(255) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(255) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(255);
OutputSelectOut(256) <= InputSelectOut(128) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(1) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(256) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(256) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(256) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(256) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(256) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(256) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(256);
OutputSelectOut(257) <= InputSelectOut(384) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(257) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(384) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(320) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(288) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(272) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(264) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(260) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(258);
OutputSelectOut(258) <= InputSelectOut(129) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(3) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(258) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(258) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(258) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(258) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(258) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(258) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(257);
OutputSelectOut(259) <= InputSelectOut(385) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(259) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(386) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(322) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(290) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(274) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(266) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(262) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(259);
OutputSelectOut(260) <= InputSelectOut(130) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(5) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(260) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(260) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(260) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(260) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(260) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(257) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(260);
OutputSelectOut(261) <= InputSelectOut(386) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(261) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(388) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(324) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(292) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(276) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(268) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(261) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(262);
OutputSelectOut(262) <= InputSelectOut(131) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(7) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(262) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(262) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(262) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(262) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(262) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(259) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(261);
OutputSelectOut(263) <= InputSelectOut(387) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(263) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(390) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(326) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(294) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(278) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(270) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(263) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(263);
OutputSelectOut(264) <= InputSelectOut(132) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(9) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(264) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(264) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(264) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(264) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(257) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(264) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(264);
OutputSelectOut(265) <= InputSelectOut(388) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(265) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(392) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(328) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(296) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(280) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(265) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(268) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(266);
OutputSelectOut(266) <= InputSelectOut(133) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(11) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(266) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(266) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(266) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(266) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(259) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(266) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(265);
OutputSelectOut(267) <= InputSelectOut(389) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(267) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(394) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(330) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(298) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(282) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(267) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(270) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(267);
OutputSelectOut(268) <= InputSelectOut(134) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(13) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(268) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(268) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(268) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(268) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(261) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(265) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(268);
OutputSelectOut(269) <= InputSelectOut(390) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(269) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(396) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(332) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(300) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(284) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(269) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(269) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(270);
OutputSelectOut(270) <= InputSelectOut(135) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(15) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(270) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(270) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(270) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(270) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(263) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(267) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(269);
OutputSelectOut(271) <= InputSelectOut(391) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(271) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(398) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(334) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(302) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(286) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(271) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(271) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(271);
OutputSelectOut(272) <= InputSelectOut(136) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(17) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(272) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(272) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(272) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(257) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(272) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(272) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(272);
OutputSelectOut(273) <= InputSelectOut(392) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(273) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(400) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(336) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(304) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(273) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(280) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(276) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(274);
OutputSelectOut(274) <= InputSelectOut(137) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(19) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(274) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(274) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(274) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(259) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(274) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(274) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(273);
OutputSelectOut(275) <= InputSelectOut(393) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(275) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(402) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(338) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(306) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(275) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(282) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(278) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(275);
OutputSelectOut(276) <= InputSelectOut(138) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(21) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(276) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(276) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(276) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(261) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(276) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(273) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(276);
OutputSelectOut(277) <= InputSelectOut(394) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(277) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(404) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(340) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(308) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(277) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(284) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(277) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(278);
OutputSelectOut(278) <= InputSelectOut(139) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(23) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(278) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(278) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(278) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(263) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(278) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(275) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(277);
OutputSelectOut(279) <= InputSelectOut(395) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(279) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(406) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(342) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(310) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(279) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(286) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(279) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(279);
OutputSelectOut(280) <= InputSelectOut(140) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(25) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(280) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(280) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(280) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(265) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(273) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(280) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(280);
OutputSelectOut(281) <= InputSelectOut(396) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(281) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(408) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(344) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(312) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(281) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(281) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(284) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(282);
OutputSelectOut(282) <= InputSelectOut(141) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(27) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(282) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(282) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(282) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(267) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(275) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(282) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(281);
OutputSelectOut(283) <= InputSelectOut(397) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(283) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(410) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(346) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(314) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(283) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(283) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(286) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(283);
OutputSelectOut(284) <= InputSelectOut(142) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(29) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(284) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(284) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(284) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(269) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(277) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(281) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(284);
OutputSelectOut(285) <= InputSelectOut(398) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(285) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(412) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(348) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(316) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(285) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(285) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(285) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(286);
OutputSelectOut(286) <= InputSelectOut(143) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(31) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(286) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(286) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(286) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(271) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(279) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(283) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(285);
OutputSelectOut(287) <= InputSelectOut(399) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(287) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(414) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(350) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(318) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(287) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(287) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(287) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(287);
OutputSelectOut(288) <= InputSelectOut(144) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(33) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(288) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(288) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(257) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(288) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(288) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(288) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(288);
OutputSelectOut(289) <= InputSelectOut(400) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(289) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(416) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(352) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(289) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(304) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(296) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(292) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(290);
OutputSelectOut(290) <= InputSelectOut(145) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(35) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(290) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(290) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(259) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(290) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(290) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(290) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(289);
OutputSelectOut(291) <= InputSelectOut(401) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(291) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(418) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(354) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(291) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(306) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(298) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(294) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(291);
OutputSelectOut(292) <= InputSelectOut(146) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(37) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(292) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(292) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(261) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(292) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(292) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(289) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(292);
OutputSelectOut(293) <= InputSelectOut(402) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(293) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(420) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(356) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(293) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(308) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(300) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(293) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(294);
OutputSelectOut(294) <= InputSelectOut(147) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(39) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(294) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(294) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(263) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(294) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(294) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(291) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(293);
OutputSelectOut(295) <= InputSelectOut(403) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(295) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(422) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(358) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(295) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(310) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(302) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(295) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(295);
OutputSelectOut(296) <= InputSelectOut(148) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(41) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(296) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(296) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(265) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(296) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(289) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(296) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(296);
OutputSelectOut(297) <= InputSelectOut(404) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(297) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(424) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(360) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(297) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(312) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(297) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(300) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(298);
OutputSelectOut(298) <= InputSelectOut(149) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(43) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(298) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(298) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(267) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(298) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(291) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(298) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(297);
OutputSelectOut(299) <= InputSelectOut(405) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(299) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(426) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(362) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(299) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(314) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(299) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(302) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(299);
OutputSelectOut(300) <= InputSelectOut(150) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(45) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(300) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(300) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(269) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(300) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(293) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(297) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(300);
OutputSelectOut(301) <= InputSelectOut(406) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(301) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(428) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(364) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(301) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(316) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(301) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(301) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(302);
OutputSelectOut(302) <= InputSelectOut(151) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(47) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(302) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(302) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(271) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(302) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(295) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(299) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(301);
OutputSelectOut(303) <= InputSelectOut(407) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(303) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(430) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(366) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(303) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(318) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(303) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(303) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(303);
OutputSelectOut(304) <= InputSelectOut(152) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(49) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(304) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(304) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(273) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(289) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(304) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(304) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(304);
OutputSelectOut(305) <= InputSelectOut(408) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(305) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(432) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(368) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(305) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(305) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(312) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(308) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(306);
OutputSelectOut(306) <= InputSelectOut(153) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(51) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(306) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(306) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(275) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(291) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(306) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(306) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(305);
OutputSelectOut(307) <= InputSelectOut(409) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(307) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(434) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(370) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(307) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(307) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(314) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(310) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(307);
OutputSelectOut(308) <= InputSelectOut(154) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(53) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(308) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(308) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(277) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(293) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(308) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(305) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(308);
OutputSelectOut(309) <= InputSelectOut(410) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(309) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(436) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(372) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(309) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(309) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(316) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(309) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(310);
OutputSelectOut(310) <= InputSelectOut(155) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(55) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(310) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(310) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(279) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(295) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(310) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(307) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(309);
OutputSelectOut(311) <= InputSelectOut(411) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(311) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(438) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(374) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(311) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(311) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(318) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(311) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(311);
OutputSelectOut(312) <= InputSelectOut(156) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(57) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(312) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(312) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(281) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(297) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(305) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(312) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(312);
OutputSelectOut(313) <= InputSelectOut(412) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(313) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(440) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(376) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(313) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(313) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(313) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(316) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(314);
OutputSelectOut(314) <= InputSelectOut(157) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(59) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(314) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(314) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(283) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(299) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(307) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(314) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(313);
OutputSelectOut(315) <= InputSelectOut(413) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(315) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(442) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(378) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(315) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(315) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(315) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(318) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(315);
OutputSelectOut(316) <= InputSelectOut(158) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(61) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(316) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(316) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(285) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(301) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(309) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(313) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(316);
OutputSelectOut(317) <= InputSelectOut(414) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(317) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(444) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(380) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(317) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(317) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(317) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(317) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(318);
OutputSelectOut(318) <= InputSelectOut(159) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(63) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(318) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(318) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(287) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(303) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(311) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(315) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(317);
OutputSelectOut(319) <= InputSelectOut(415) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(319) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(446) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(382) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(319) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(319) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(319) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(319) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(319);
OutputSelectOut(320) <= InputSelectOut(160) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(65) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(320) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(257) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(320) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(320) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(320) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(320) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(320);
OutputSelectOut(321) <= InputSelectOut(416) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(321) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(448) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(321) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(352) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(336) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(328) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(324) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(322);
OutputSelectOut(322) <= InputSelectOut(161) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(67) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(322) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(259) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(322) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(322) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(322) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(322) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(321);
OutputSelectOut(323) <= InputSelectOut(417) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(323) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(450) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(323) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(354) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(338) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(330) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(326) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(323);
OutputSelectOut(324) <= InputSelectOut(162) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(69) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(324) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(261) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(324) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(324) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(324) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(321) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(324);
OutputSelectOut(325) <= InputSelectOut(418) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(325) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(452) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(325) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(356) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(340) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(332) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(325) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(326);
OutputSelectOut(326) <= InputSelectOut(163) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(71) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(326) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(263) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(326) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(326) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(326) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(323) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(325);
OutputSelectOut(327) <= InputSelectOut(419) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(327) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(454) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(327) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(358) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(342) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(334) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(327) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(327);
OutputSelectOut(328) <= InputSelectOut(164) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(73) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(328) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(265) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(328) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(328) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(321) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(328) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(328);
OutputSelectOut(329) <= InputSelectOut(420) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(329) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(456) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(329) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(360) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(344) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(329) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(332) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(330);
OutputSelectOut(330) <= InputSelectOut(165) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(75) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(330) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(267) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(330) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(330) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(323) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(330) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(329);
OutputSelectOut(331) <= InputSelectOut(421) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(331) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(458) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(331) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(362) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(346) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(331) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(334) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(331);
OutputSelectOut(332) <= InputSelectOut(166) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(77) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(332) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(269) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(332) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(332) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(325) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(329) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(332);
OutputSelectOut(333) <= InputSelectOut(422) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(333) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(460) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(333) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(364) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(348) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(333) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(333) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(334);
OutputSelectOut(334) <= InputSelectOut(167) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(79) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(334) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(271) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(334) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(334) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(327) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(331) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(333);
OutputSelectOut(335) <= InputSelectOut(423) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(335) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(462) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(335) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(366) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(350) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(335) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(335) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(335);
OutputSelectOut(336) <= InputSelectOut(168) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(81) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(336) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(273) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(336) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(321) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(336) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(336) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(336);
OutputSelectOut(337) <= InputSelectOut(424) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(337) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(464) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(337) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(368) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(337) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(344) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(340) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(338);
OutputSelectOut(338) <= InputSelectOut(169) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(83) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(338) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(275) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(338) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(323) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(338) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(338) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(337);
OutputSelectOut(339) <= InputSelectOut(425) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(339) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(466) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(339) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(370) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(339) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(346) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(342) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(339);
OutputSelectOut(340) <= InputSelectOut(170) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(85) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(340) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(277) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(340) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(325) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(340) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(337) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(340);
OutputSelectOut(341) <= InputSelectOut(426) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(341) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(468) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(341) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(372) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(341) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(348) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(341) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(342);
OutputSelectOut(342) <= InputSelectOut(171) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(87) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(342) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(279) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(342) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(327) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(342) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(339) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(341);
OutputSelectOut(343) <= InputSelectOut(427) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(343) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(470) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(343) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(374) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(343) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(350) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(343) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(343);
OutputSelectOut(344) <= InputSelectOut(172) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(89) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(344) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(281) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(344) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(329) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(337) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(344) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(344);
OutputSelectOut(345) <= InputSelectOut(428) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(345) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(472) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(345) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(376) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(345) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(345) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(348) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(346);
OutputSelectOut(346) <= InputSelectOut(173) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(91) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(346) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(283) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(346) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(331) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(339) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(346) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(345);
OutputSelectOut(347) <= InputSelectOut(429) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(347) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(474) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(347) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(378) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(347) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(347) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(350) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(347);
OutputSelectOut(348) <= InputSelectOut(174) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(93) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(348) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(285) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(348) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(333) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(341) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(345) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(348);
OutputSelectOut(349) <= InputSelectOut(430) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(349) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(476) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(349) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(380) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(349) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(349) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(349) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(350);
OutputSelectOut(350) <= InputSelectOut(175) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(95) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(350) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(287) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(350) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(335) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(343) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(347) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(349);
OutputSelectOut(351) <= InputSelectOut(431) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(351) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(478) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(351) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(382) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(351) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(351) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(351) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(351);
OutputSelectOut(352) <= InputSelectOut(176) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(97) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(352) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(289) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(321) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(352) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(352) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(352) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(352);
OutputSelectOut(353) <= InputSelectOut(432) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(353) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(480) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(353) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(353) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(368) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(360) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(356) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(354);
OutputSelectOut(354) <= InputSelectOut(177) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(99) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(354) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(291) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(323) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(354) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(354) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(354) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(353);
OutputSelectOut(355) <= InputSelectOut(433) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(355) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(482) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(355) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(355) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(370) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(362) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(358) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(355);
OutputSelectOut(356) <= InputSelectOut(178) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(101) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(356) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(293) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(325) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(356) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(356) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(353) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(356);
OutputSelectOut(357) <= InputSelectOut(434) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(357) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(484) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(357) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(357) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(372) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(364) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(357) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(358);
OutputSelectOut(358) <= InputSelectOut(179) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(103) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(358) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(295) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(327) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(358) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(358) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(355) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(357);
OutputSelectOut(359) <= InputSelectOut(435) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(359) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(486) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(359) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(359) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(374) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(366) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(359) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(359);
OutputSelectOut(360) <= InputSelectOut(180) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(105) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(360) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(297) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(329) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(360) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(353) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(360) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(360);
OutputSelectOut(361) <= InputSelectOut(436) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(361) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(488) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(361) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(361) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(376) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(361) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(364) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(362);
OutputSelectOut(362) <= InputSelectOut(181) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(107) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(362) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(299) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(331) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(362) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(355) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(362) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(361);
OutputSelectOut(363) <= InputSelectOut(437) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(363) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(490) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(363) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(363) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(378) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(363) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(366) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(363);
OutputSelectOut(364) <= InputSelectOut(182) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(109) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(364) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(301) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(333) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(364) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(357) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(361) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(364);
OutputSelectOut(365) <= InputSelectOut(438) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(365) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(492) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(365) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(365) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(380) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(365) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(365) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(366);
OutputSelectOut(366) <= InputSelectOut(183) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(111) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(366) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(303) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(335) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(366) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(359) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(363) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(365);
OutputSelectOut(367) <= InputSelectOut(439) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(367) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(494) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(367) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(367) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(382) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(367) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(367) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(367);
OutputSelectOut(368) <= InputSelectOut(184) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(113) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(368) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(305) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(337) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(353) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(368) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(368) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(368);
OutputSelectOut(369) <= InputSelectOut(440) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(369) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(496) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(369) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(369) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(369) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(376) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(372) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(370);
OutputSelectOut(370) <= InputSelectOut(185) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(115) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(370) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(307) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(339) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(355) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(370) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(370) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(369);
OutputSelectOut(371) <= InputSelectOut(441) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(371) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(498) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(371) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(371) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(371) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(378) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(374) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(371);
OutputSelectOut(372) <= InputSelectOut(186) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(117) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(372) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(309) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(341) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(357) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(372) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(369) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(372);
OutputSelectOut(373) <= InputSelectOut(442) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(373) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(500) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(373) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(373) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(373) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(380) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(373) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(374);
OutputSelectOut(374) <= InputSelectOut(187) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(119) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(374) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(311) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(343) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(359) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(374) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(371) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(373);
OutputSelectOut(375) <= InputSelectOut(443) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(375) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(502) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(375) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(375) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(375) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(382) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(375) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(375);
OutputSelectOut(376) <= InputSelectOut(188) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(121) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(376) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(313) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(345) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(361) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(369) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(376) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(376);
OutputSelectOut(377) <= InputSelectOut(444) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(377) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(504) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(377) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(377) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(377) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(377) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(380) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(378);
OutputSelectOut(378) <= InputSelectOut(189) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(123) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(378) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(315) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(347) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(363) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(371) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(378) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(377);
OutputSelectOut(379) <= InputSelectOut(445) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(379) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(506) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(379) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(379) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(379) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(379) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(382) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(379);
OutputSelectOut(380) <= InputSelectOut(190) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(125) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(380) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(317) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(349) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(365) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(373) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(377) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(380);
OutputSelectOut(381) <= InputSelectOut(446) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(381) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(508) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(381) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(381) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(381) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(381) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(381) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(382);
OutputSelectOut(382) <= InputSelectOut(191) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(127) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(382) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(319) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(351) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(367) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(375) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(379) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(381);
OutputSelectOut(383) <= InputSelectOut(447) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(383) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(510) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(383) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(383) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(383) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(383) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(383) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(383);
OutputSelectOut(384) <= InputSelectOut(192) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(129) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(257) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(384) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(384) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(384) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(384) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(384) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(384);
OutputSelectOut(385) <= InputSelectOut(448) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(385) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(385) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(448) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(416) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(400) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(392) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(388) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(386);
OutputSelectOut(386) <= InputSelectOut(193) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(131) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(259) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(386) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(386) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(386) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(386) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(386) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(385);
OutputSelectOut(387) <= InputSelectOut(449) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(387) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(387) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(450) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(418) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(402) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(394) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(390) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(387);
OutputSelectOut(388) <= InputSelectOut(194) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(133) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(261) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(388) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(388) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(388) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(388) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(385) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(388);
OutputSelectOut(389) <= InputSelectOut(450) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(389) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(389) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(452) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(420) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(404) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(396) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(389) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(390);
OutputSelectOut(390) <= InputSelectOut(195) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(135) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(263) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(390) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(390) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(390) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(390) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(387) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(389);
OutputSelectOut(391) <= InputSelectOut(451) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(391) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(391) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(454) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(422) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(406) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(398) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(391) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(391);
OutputSelectOut(392) <= InputSelectOut(196) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(137) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(265) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(392) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(392) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(392) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(385) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(392) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(392);
OutputSelectOut(393) <= InputSelectOut(452) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(393) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(393) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(456) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(424) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(408) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(393) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(396) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(394);
OutputSelectOut(394) <= InputSelectOut(197) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(139) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(267) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(394) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(394) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(394) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(387) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(394) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(393);
OutputSelectOut(395) <= InputSelectOut(453) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(395) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(395) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(458) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(426) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(410) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(395) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(398) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(395);
OutputSelectOut(396) <= InputSelectOut(198) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(141) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(269) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(396) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(396) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(396) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(389) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(393) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(396);
OutputSelectOut(397) <= InputSelectOut(454) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(397) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(397) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(460) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(428) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(412) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(397) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(397) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(398);
OutputSelectOut(398) <= InputSelectOut(199) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(143) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(271) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(398) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(398) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(398) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(391) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(395) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(397);
OutputSelectOut(399) <= InputSelectOut(455) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(399) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(399) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(462) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(430) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(414) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(399) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(399) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(399);
OutputSelectOut(400) <= InputSelectOut(200) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(145) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(273) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(400) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(400) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(385) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(400) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(400) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(400);
OutputSelectOut(401) <= InputSelectOut(456) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(401) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(401) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(464) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(432) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(401) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(408) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(404) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(402);
OutputSelectOut(402) <= InputSelectOut(201) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(147) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(275) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(402) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(402) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(387) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(402) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(402) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(401);
OutputSelectOut(403) <= InputSelectOut(457) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(403) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(403) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(466) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(434) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(403) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(410) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(406) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(403);
OutputSelectOut(404) <= InputSelectOut(202) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(149) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(277) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(404) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(404) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(389) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(404) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(401) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(404);
OutputSelectOut(405) <= InputSelectOut(458) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(405) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(405) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(468) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(436) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(405) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(412) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(405) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(406);
OutputSelectOut(406) <= InputSelectOut(203) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(151) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(279) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(406) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(406) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(391) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(406) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(403) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(405);
OutputSelectOut(407) <= InputSelectOut(459) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(407) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(407) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(470) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(438) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(407) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(414) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(407) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(407);
OutputSelectOut(408) <= InputSelectOut(204) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(153) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(281) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(408) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(408) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(393) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(401) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(408) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(408);
OutputSelectOut(409) <= InputSelectOut(460) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(409) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(409) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(472) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(440) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(409) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(409) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(412) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(410);
OutputSelectOut(410) <= InputSelectOut(205) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(155) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(283) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(410) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(410) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(395) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(403) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(410) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(409);
OutputSelectOut(411) <= InputSelectOut(461) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(411) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(411) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(474) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(442) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(411) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(411) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(414) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(411);
OutputSelectOut(412) <= InputSelectOut(206) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(157) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(285) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(412) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(412) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(397) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(405) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(409) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(412);
OutputSelectOut(413) <= InputSelectOut(462) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(413) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(413) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(476) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(444) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(413) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(413) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(413) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(414);
OutputSelectOut(414) <= InputSelectOut(207) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(159) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(287) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(414) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(414) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(399) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(407) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(411) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(413);
OutputSelectOut(415) <= InputSelectOut(463) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(415) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(415) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(478) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(446) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(415) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(415) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(415) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(415);
OutputSelectOut(416) <= InputSelectOut(208) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(161) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(289) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(416) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(385) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(416) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(416) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(416) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(416);
OutputSelectOut(417) <= InputSelectOut(464) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(417) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(417) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(480) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(417) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(432) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(424) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(420) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(418);
OutputSelectOut(418) <= InputSelectOut(209) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(163) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(291) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(418) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(387) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(418) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(418) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(418) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(417);
OutputSelectOut(419) <= InputSelectOut(465) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(419) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(419) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(482) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(419) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(434) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(426) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(422) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(419);
OutputSelectOut(420) <= InputSelectOut(210) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(165) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(293) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(420) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(389) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(420) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(420) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(417) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(420);
OutputSelectOut(421) <= InputSelectOut(466) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(421) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(421) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(484) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(421) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(436) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(428) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(421) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(422);
OutputSelectOut(422) <= InputSelectOut(211) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(167) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(295) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(422) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(391) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(422) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(422) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(419) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(421);
OutputSelectOut(423) <= InputSelectOut(467) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(423) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(423) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(486) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(423) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(438) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(430) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(423) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(423);
OutputSelectOut(424) <= InputSelectOut(212) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(169) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(297) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(424) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(393) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(424) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(417) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(424) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(424);
OutputSelectOut(425) <= InputSelectOut(468) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(425) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(425) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(488) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(425) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(440) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(425) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(428) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(426);
OutputSelectOut(426) <= InputSelectOut(213) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(171) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(299) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(426) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(395) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(426) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(419) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(426) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(425);
OutputSelectOut(427) <= InputSelectOut(469) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(427) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(427) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(490) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(427) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(442) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(427) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(430) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(427);
OutputSelectOut(428) <= InputSelectOut(214) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(173) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(301) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(428) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(397) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(428) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(421) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(425) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(428);
OutputSelectOut(429) <= InputSelectOut(470) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(429) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(429) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(492) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(429) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(444) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(429) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(429) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(430);
OutputSelectOut(430) <= InputSelectOut(215) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(175) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(303) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(430) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(399) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(430) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(423) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(427) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(429);
OutputSelectOut(431) <= InputSelectOut(471) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(431) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(431) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(494) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(431) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(446) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(431) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(431) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(431);
OutputSelectOut(432) <= InputSelectOut(216) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(177) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(305) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(432) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(401) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(417) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(432) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(432) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(432);
OutputSelectOut(433) <= InputSelectOut(472) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(433) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(433) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(496) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(433) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(433) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(440) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(436) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(434);
OutputSelectOut(434) <= InputSelectOut(217) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(179) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(307) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(434) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(403) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(419) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(434) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(434) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(433);
OutputSelectOut(435) <= InputSelectOut(473) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(435) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(435) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(498) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(435) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(435) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(442) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(438) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(435);
OutputSelectOut(436) <= InputSelectOut(218) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(181) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(309) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(436) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(405) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(421) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(436) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(433) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(436);
OutputSelectOut(437) <= InputSelectOut(474) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(437) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(437) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(500) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(437) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(437) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(444) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(437) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(438);
OutputSelectOut(438) <= InputSelectOut(219) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(183) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(311) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(438) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(407) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(423) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(438) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(435) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(437);
OutputSelectOut(439) <= InputSelectOut(475) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(439) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(439) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(502) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(439) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(439) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(446) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(439) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(439);
OutputSelectOut(440) <= InputSelectOut(220) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(185) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(313) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(440) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(409) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(425) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(433) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(440) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(440);
OutputSelectOut(441) <= InputSelectOut(476) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(441) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(441) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(504) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(441) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(441) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(441) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(444) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(442);
OutputSelectOut(442) <= InputSelectOut(221) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(187) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(315) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(442) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(411) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(427) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(435) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(442) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(441);
OutputSelectOut(443) <= InputSelectOut(477) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(443) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(443) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(506) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(443) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(443) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(443) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(446) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(443);
OutputSelectOut(444) <= InputSelectOut(222) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(189) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(317) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(444) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(413) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(429) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(437) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(441) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(444);
OutputSelectOut(445) <= InputSelectOut(478) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(445) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(445) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(508) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(445) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(445) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(445) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(445) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(446);
OutputSelectOut(446) <= InputSelectOut(223) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(191) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(319) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(446) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(415) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(431) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(439) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(443) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(445);
OutputSelectOut(447) <= InputSelectOut(479) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(447) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(447) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(510) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(447) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(447) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(447) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(447) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(447);
OutputSelectOut(448) <= InputSelectOut(224) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(193) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(321) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(385) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(448) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(448) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(448) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(448) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(448);
OutputSelectOut(449) <= InputSelectOut(480) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(449) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(449) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(449) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(480) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(464) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(456) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(452) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(450);
OutputSelectOut(450) <= InputSelectOut(225) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(195) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(323) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(387) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(450) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(450) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(450) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(450) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(449);
OutputSelectOut(451) <= InputSelectOut(481) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(451) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(451) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(451) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(482) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(466) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(458) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(454) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(451);
OutputSelectOut(452) <= InputSelectOut(226) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(197) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(325) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(389) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(452) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(452) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(452) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(449) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(452);
OutputSelectOut(453) <= InputSelectOut(482) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(453) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(453) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(453) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(484) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(468) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(460) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(453) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(454);
OutputSelectOut(454) <= InputSelectOut(227) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(199) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(327) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(391) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(454) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(454) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(454) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(451) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(453);
OutputSelectOut(455) <= InputSelectOut(483) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(455) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(455) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(455) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(486) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(470) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(462) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(455) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(455);
OutputSelectOut(456) <= InputSelectOut(228) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(201) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(329) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(393) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(456) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(456) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(449) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(456) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(456);
OutputSelectOut(457) <= InputSelectOut(484) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(457) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(457) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(457) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(488) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(472) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(457) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(460) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(458);
OutputSelectOut(458) <= InputSelectOut(229) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(203) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(331) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(395) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(458) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(458) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(451) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(458) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(457);
OutputSelectOut(459) <= InputSelectOut(485) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(459) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(459) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(459) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(490) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(474) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(459) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(462) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(459);
OutputSelectOut(460) <= InputSelectOut(230) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(205) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(333) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(397) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(460) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(460) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(453) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(457) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(460);
OutputSelectOut(461) <= InputSelectOut(486) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(461) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(461) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(461) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(492) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(476) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(461) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(461) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(462);
OutputSelectOut(462) <= InputSelectOut(231) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(207) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(335) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(399) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(462) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(462) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(455) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(459) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(461);
OutputSelectOut(463) <= InputSelectOut(487) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(463) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(463) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(463) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(494) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(478) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(463) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(463) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(463);
OutputSelectOut(464) <= InputSelectOut(232) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(209) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(337) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(401) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(464) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(449) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(464) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(464) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(464);
OutputSelectOut(465) <= InputSelectOut(488) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(465) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(465) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(465) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(496) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(465) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(472) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(468) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(466);
OutputSelectOut(466) <= InputSelectOut(233) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(211) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(339) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(403) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(466) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(451) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(466) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(466) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(465);
OutputSelectOut(467) <= InputSelectOut(489) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(467) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(467) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(467) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(498) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(467) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(474) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(470) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(467);
OutputSelectOut(468) <= InputSelectOut(234) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(213) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(341) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(405) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(468) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(453) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(468) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(465) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(468);
OutputSelectOut(469) <= InputSelectOut(490) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(469) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(469) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(469) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(500) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(469) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(476) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(469) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(470);
OutputSelectOut(470) <= InputSelectOut(235) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(215) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(343) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(407) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(470) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(455) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(470) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(467) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(469);
OutputSelectOut(471) <= InputSelectOut(491) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(471) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(471) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(471) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(502) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(471) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(478) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(471) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(471);
OutputSelectOut(472) <= InputSelectOut(236) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(217) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(345) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(409) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(472) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(457) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(465) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(472) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(472);
OutputSelectOut(473) <= InputSelectOut(492) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(473) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(473) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(473) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(504) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(473) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(473) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(476) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(474);
OutputSelectOut(474) <= InputSelectOut(237) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(219) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(347) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(411) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(474) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(459) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(467) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(474) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(473);
OutputSelectOut(475) <= InputSelectOut(493) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(475) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(475) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(475) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(506) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(475) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(475) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(478) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(475);
OutputSelectOut(476) <= InputSelectOut(238) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(221) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(349) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(413) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(476) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(461) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(469) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(473) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(476);
OutputSelectOut(477) <= InputSelectOut(494) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(477) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(477) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(477) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(508) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(477) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(477) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(477) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(478);
OutputSelectOut(478) <= InputSelectOut(239) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(223) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(351) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(415) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(478) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(463) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(471) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(475) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(477);
OutputSelectOut(479) <= InputSelectOut(495) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(479) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(479) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(479) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(510) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(479) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(479) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(479) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(479);
OutputSelectOut(480) <= InputSelectOut(240) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(225) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(353) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(417) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(449) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(480) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(480) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(480) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(480);
OutputSelectOut(481) <= InputSelectOut(496) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(481) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(481) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(481) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(481) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(496) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(488) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(484) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(482);
OutputSelectOut(482) <= InputSelectOut(241) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(227) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(355) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(419) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(451) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(482) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(482) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(482) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(481);
OutputSelectOut(483) <= InputSelectOut(497) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(483) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(483) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(483) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(483) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(498) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(490) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(486) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(483);
OutputSelectOut(484) <= InputSelectOut(242) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(229) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(357) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(421) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(453) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(484) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(484) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(481) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(484);
OutputSelectOut(485) <= InputSelectOut(498) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(485) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(485) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(485) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(485) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(500) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(492) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(485) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(486);
OutputSelectOut(486) <= InputSelectOut(243) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(231) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(359) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(423) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(455) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(486) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(486) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(483) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(485);
OutputSelectOut(487) <= InputSelectOut(499) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(487) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(487) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(487) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(487) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(502) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(494) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(487) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(487);
OutputSelectOut(488) <= InputSelectOut(244) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(233) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(361) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(425) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(457) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(488) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(481) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(488) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(488);
OutputSelectOut(489) <= InputSelectOut(500) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(489) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(489) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(489) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(489) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(504) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(489) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(492) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(490);
OutputSelectOut(490) <= InputSelectOut(245) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(235) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(363) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(427) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(459) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(490) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(483) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(490) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(489);
OutputSelectOut(491) <= InputSelectOut(501) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(491) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(491) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(491) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(491) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(506) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(491) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(494) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(491);
OutputSelectOut(492) <= InputSelectOut(246) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(237) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(365) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(429) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(461) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(492) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(485) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(489) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(492);
OutputSelectOut(493) <= InputSelectOut(502) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(493) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(493) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(493) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(493) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(508) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(493) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(493) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(494);
OutputSelectOut(494) <= InputSelectOut(247) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(239) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(367) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(431) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(463) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(494) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(487) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(491) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(493);
OutputSelectOut(495) <= InputSelectOut(503) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(495) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(495) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(495) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(495) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(510) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(495) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(495) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(495);
OutputSelectOut(496) <= InputSelectOut(248) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(241) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(369) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(433) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(465) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(481) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(496) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(496) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(496);
OutputSelectOut(497) <= InputSelectOut(504) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(497) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(497) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(497) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(497) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(497) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(504) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(500) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(498);
OutputSelectOut(498) <= InputSelectOut(249) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(243) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(371) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(435) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(467) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(483) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(498) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(498) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(497);
OutputSelectOut(499) <= InputSelectOut(505) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(499) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(499) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(499) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(499) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(499) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(506) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(502) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(499);
OutputSelectOut(500) <= InputSelectOut(250) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(245) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(373) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(437) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(469) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(485) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(500) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(497) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(500);
OutputSelectOut(501) <= InputSelectOut(506) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(501) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(501) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(501) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(501) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(501) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(508) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(501) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(502);
OutputSelectOut(502) <= InputSelectOut(251) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(247) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(375) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(439) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(471) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(487) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(502) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(499) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(501);
OutputSelectOut(503) <= InputSelectOut(507) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(503) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(503) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(503) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(503) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(503) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(510) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(503) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(503);
OutputSelectOut(504) <= InputSelectOut(252) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(249) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(377) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(441) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(473) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(489) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(497) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(504) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(504);
OutputSelectOut(505) <= InputSelectOut(508) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(505) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(505) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(505) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(505) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(505) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(505) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(508) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(506);
OutputSelectOut(506) <= InputSelectOut(253) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(251) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(379) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(443) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(475) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(491) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(499) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(506) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(505);
OutputSelectOut(507) <= InputSelectOut(509) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(507) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(507) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(507) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(507) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(507) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(507) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(510) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(507);
OutputSelectOut(508) <= InputSelectOut(254) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(253) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(381) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(445) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(477) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(493) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(501) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(505) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(508);
OutputSelectOut(509) <= InputSelectOut(510) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(509) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(509) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(509) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(509) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(509) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(509) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(509) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(510);
OutputSelectOut(510) <= InputSelectOut(255) WHEN ControlSelectOut = "0000" ELSE
			 InputSelectOut(255) WHEN ControlSelectOut = "0001" ELSE
			 InputSelectOut(383) WHEN ControlSelectOut = "0010" ELSE
			 InputSelectOut(447) WHEN ControlSelectOut = "0011" ELSE
			 InputSelectOut(479) WHEN ControlSelectOut = "0100" ELSE
			 InputSelectOut(495) WHEN ControlSelectOut = "0101" ELSE
			 InputSelectOut(503) WHEN ControlSelectOut = "0110" ELSE
			 InputSelectOut(507) WHEN ControlSelectOut = "0111" ELSE
			 InputSelectOut(509);
OutputSelectOut(511) <= InputSelectOut(511);


END Behavioral;