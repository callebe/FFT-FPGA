library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT1024p_4 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT1024p_4;

architecture Behavioral of ROMFFT1024p_4 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 5 
	constant ROM_tb : ROM := (
		0 => "011000000110111110101",
		1 => "011000000110111110101",
		2 => "011000000110111110101",
		3 => "011011101110001010000",
		4 => "011011101110001010000",
		5 => "011011101110001010000",
		6 => "011100000100001010011",
		7 => "011100000100001010011",
		8 => "011100000100001010011",
		9 => "001010011100001010111",
		10 => "001010011100001010111",
		11 => "001010011100001010111",
		12 => "011010100100001010010",
		13 => "011010100100001010010",
		14 => "011010100100001010010",
		15 => "001001100101101110000",
		16 => "001001100101101110000",
		17 => "001001100101101110000",
		18 => "001001011100001010101",
		19 => "001001011100001010101",
		20 => "001001011100001010101",
		21 => "011010100100001010010",
		22 => "011010100100001010010",
		23 => "011010100100001010010",
		24 => "001000111100001110011",
		25 => "001000111100001110011",
		26 => "001000111100001110011",
		27 => "011000001101100010011",
		28 => "011000001101100010011",
		29 => "011000001101100010011",
		30 => "011000000101111011000",
		31 => "011000000101111011000",
		32 => "011000000101111011000",
		33 => "001001011100001010100",
		34 => "001001011100001010100",
		35 => "001001011100001010100",
		36 => "011001111100011110010",
		37 => "011001111100011110010",
		38 => "011001111100011110010",
		39 => "011000001100101010110",
		40 => "011000001100101010110",
		41 => "011000001100101010110",
		42 => "001010011100011110010",
		43 => "001010011100011110010",
		44 => "001010011100011110010",
		45 => "011000011100111010000",
		46 => "011000011100111010000",
		47 => "011000011100111010000",
		48 => "011001100100001110000",
		49 => "011001100100001110000",
		50 => "011001100100001110000",
		51 => "011000101100101010100",
		52 => "011000101100101010100",
		53 => "011000101100101010100",
		54 => "001011011100001110010",
		55 => "001011011100001110010",
		56 => "001011011100001110010",
		57 => "001001111100011110010",
		58 => "001001111100011110010",
		59 => "001001111100011110010",
		60 => "011000000101001010010",
		61 => "011000000101001010010",
		62 => "011000000101001010010",
		63 => "011000000100111010001",
		64 => "011000000100111010001",
		65 => "011000000100111010001",
		66 => "011000001101100010011",
		67 => "011000001101100010011",
		68 => "011000001101100010011",
		69 => "001000110100001010011",
		70 => "001000110100001010011",
		71 => "001000110100001010011",
		72 => "011010100100001110010",
		73 => "011010100100001110010",
		74 => "011010100100001110010",
		75 => "011000000101011010010",
		76 => "011000000101011010010",
		77 => "011000000101011010010",
		78 => "011000000101101010011",
		79 => "011000000101101010011",
		80 => "011000000101101010011",
		81 => "011000000101011010010",
		82 => "011000000101011010010",
		83 => "011000000101011010010",
		84 => "011000000101111010100",
		85 => "011000000101111010100",
		86 => "011000000101111010100",
		87 => "001001111110001010000",
		88 => "001001111110001010000",
		89 => "001001111110001010000",
		90 => "011000011110001010110",
		91 => "011000011110001010110",
		92 => "011000011110001010110",
		93 => "011000000110111010101",
		94 => "011000000110111010101",
		95 => "011000000110111010101",
		96 => "011000000110011110100",
		97 => "011000000110011110100",
		98 => "011000000110011110100",
		99 => "011000000101110011001",
		100 => "011000000101110011001",
		101 => "011000000101110011001",
		102 => "011000001110100010101",
		103 => "011000001110100010101",
		104 => "011000001110100010101",
		105 => "001001111100001010101",
		106 => "001001111100001010101",
		107 => "001001111100001010101",
		108 => "011000000100111010110",
		109 => "011000000100111010110",
		110 => "011000000100111010110",
		111 => "001011011100001010111",
		112 => "001011011100001010111",
		113 => "001011011100001010111",
		114 => "001001111100001010110",
		115 => "001001111100001010110",
		116 => "001001111100001010110",
		117 => "011001011100111010000",
		118 => "011001011100111010000",
		119 => "011001011100111010000",
		120 => "011001011100001010011",
		121 => "011001011100001010011",
		122 => "011001011100001010011",
		123 => "011000000101101010011",
		124 => "011000000101101010011",
		125 => "011000000101101010011",
		126 => "011000111100001010011",
		127 => "011000111100001010011",
		128 => "011000111100001010011",
		129 => "011000001101110010011",
		130 => "011000001101110010011",
		131 => "011000001101110010011",
		132 => "011000000101011010011",
		133 => "011000000101011010011",
		134 => "011000000101011010011",
		135 => "011000001110100010101",
		136 => "011000001110100010101",
		137 => "011000001110100010101",
		138 => "011000010100111010110",
		139 => "011000010100111010110",
		140 => "011000010100111010110",
		141 => "011000000110011010100",
		142 => "011000000110011010100",
		143 => "011000000110011010100",
		144 => "001010011100001011001",
		145 => "001010011100001011001",
		146 => "001010011100001011001",
		147 => "011000000101110011001",
		148 => "011000000101110011001",
		149 => "011000000101110011001",
		150 => "011000001110100010101",
		151 => "011000001110100010101",
		152 => "011000001110100010101",
		153 => "001000011101011010010",
		154 => "001000011101011010010",
		155 => "001000011101011010010",
		156 => "011000001101110010011",
		157 => "011000001101110010011",
		158 => "011000001101110010011",
		159 => "011000111100111010000",
		160 => "011000111100111010000",
		161 => "011000111100111010000",
		162 => "011011000100001010011",
		163 => "011011000100001010011",
		164 => "011011000100001010011",
		165 => "011001100100001010010",
		166 => "011001100100001010010",
		167 => "011001100100001010010",
		168 => "011001100100001110010",
		169 => "011001100100001110010",
		170 => "011001100100001110010",
		171 => "011000000101101010011",
		172 => "011000000101101010011",
		173 => "011000000101101010011",
		174 => "011001100100001110001",
		175 => "011001100100001110001",
		176 => "011001100100001110001",
		177 => "011000001101110010011",
		178 => "011000001101110010011",
		179 => "011000001101110010011",
		180 => "011010100100001110011",
		181 => "011010100100001110011",
		182 => "011010100100001110011",
		183 => "011000001110100010101",
		184 => "011000001110100010101",
		185 => "011000001110100010101",
		186 => "011000000101110011001",
		187 => "011000000101110011001",
		188 => "011000000101110011001",
		189 => "001010011110011010000",
		190 => "001010011110011010000",
		191 => "001010011110011010000",
		192 => "011000000101111110011",
		193 => "011000000101111110011",
		194 => "011000000101111110011",
		195 => "001010111100001010101",
		196 => "001010111100001010101",
		197 => "001010111100001010101",
		198 => "011001011101001010000",
		199 => "011001011101001010000",
		200 => "011001011101001010000",
		201 => "001000111100011110011",
		202 => "001000111100011110011",
		203 => "001000111100011110011",
		204 => "011000101100111010001",
		205 => "011000101100111010001",
		206 => "011000101100111010001",
		207 => "011001011100001010100",
		208 => "011001011100001010100",
		209 => "011001011100001010100",
		210 => "011000000101011010101",
		211 => "011000000101011010101",
		212 => "011000000101011010101",
		213 => "011011100100001110011",
		214 => "011011100100001110011",
		215 => "011011100100001110011",
		216 => "001001111100001010111",
		217 => "001001111100001010111",
		218 => "001001111100001010111",
		219 => "011010100100001010101",
		220 => "011010100100001010101",
		221 => "011010100100001010101",
		222 => "011010000100001010010",
		223 => "011010000100001010010",
		224 => "011010000100001010010",
		225 => "001000100100111010001",
		226 => "001000100100111010001",
		227 => "001000100100111010001",
		228 => "001000000100101110110",
		229 => "001000000100101110110",
		230 => "001000000100101110110",
		231 => "011010000100001110010",
		232 => "011010000100001110010",
		233 => "011010000100001110010",
		234 => "011000000101011010101",
		235 => "011000000101011010101",
		236 => "011000000101011010101",
		237 => "011000000101111010011",
		238 => "011000000101111010011",
		239 => "011000000101111010011",
		240 => "011000000101111110011",
		241 => "011000000101111110011",
		242 => "011000000101111110011",
		243 => "001010111100001010101",
		244 => "001010111100001010101",
		245 => "001010111100001010101",
		246 => "011001011101001010000",
		247 => "011001011101001010000",
		248 => "011001011101001010000",
		249 => "001000111100011110011",
		250 => "001000111100011110011",
		251 => "001000111100011110011",
		252 => "011000101100111010001",
		253 => "011000101100111010001",
		254 => "011000101100111010001",
		255 => "011001011100001010100",
		256 => "011001011100001010100",
		257 => "011001011100001010100",
		258 => "011000000101011010101",
		259 => "011000000101011010101",
		260 => "011000000101011010101",
		261 => "011011100100001110011",
		262 => "011011100100001110011",
		263 => "011011100100001110011",
		264 => "001001111100001010111",
		265 => "001001111100001010111",
		266 => "001001111100001010111",
		267 => "011010100100001010101",
		268 => "011010100100001010101",
		269 => "011010100100001010101",
		270 => "011010000100001010010",
		271 => "011010000100001010010",
		272 => "011010000100001010010",
		273 => "001000100100111010001",
		274 => "001000100100111010001",
		275 => "001000100100111010001",
		276 => "001000000100101110110",
		277 => "001000000100101110110",
		278 => "001000000100101110110",
		279 => "011010000100001110010",
		280 => "011010000100001110010",
		281 => "011010000100001110010",
		282 => "011000000101011010101",
		283 => "011000000101011010101",
		284 => "011000000101011010101",
		285 => "011000000101111010011",
		286 => "011000000101111010011",
		287 => "011000000101111010011",
		288 => "011010100100001110100",
		289 => "011010100100001110100",
		290 => "011010100100001110100",
		291 => "011000001101100010011",
		292 => "011000001101100010011",
		293 => "011000001101100010011",
		294 => "111011010100001010011",
		295 => "111011010100001010011",
		296 => "111011010100001010011",
		297 => "011010100100001010100",
		298 => "011010100100001010100",
		299 => "011010100100001010100",
		300 => "011010100100001110100",
		301 => "011010100100001110100",
		302 => "011010100100001110100",
		303 => "011000001101100010011",
		304 => "011000001101100010011",
		305 => "011000001101100010011",
		306 => "011000001101100010011",
		307 => "011000001101100010011",
		308 => "011000001101100010011",
		309 => "011010100100001010100",
		310 => "011010100100001010100",
		311 => "011010100100001010100",
		312 => "011010100100001110100",
		313 => "011010100100001110100",
		314 => "011010100100001110100",
		315 => "011000001101100010011",
		316 => "011000001101100010011",
		317 => "011000001101100010011",
		318 => "111011010100001010011",
		319 => "111011010100001010011",
		320 => "111011010100001010011",
		321 => "011010100100001010100",
		322 => "011010100100001010100",
		323 => "011010100100001010100",
		324 => "011010100100001110100",
		325 => "011010100100001110100",
		326 => "011010100100001110100",
		327 => "011000001101100010011",
		328 => "011000001101100010011",
		329 => "011000001101100010011",
		330 => "011000001101100010011",
		331 => "011000001101100010011",
		332 => "011000001101100010011",
		333 => "011010100100001010100",
		334 => "011010100100001010100",
		335 => "011010100100001010100",
		336 => "011010100100001110100",
		337 => "011010100100001110100",
		338 => "011010100100001110100",
		339 => "011000001101100010011",
		340 => "011000001101100010011",
		341 => "011000001101100010011",
		342 => "111011010100001010011",
		343 => "111011010100001010011",
		344 => "111011010100001010011",
		345 => "011010100100001010100",
		346 => "011010100100001010100",
		347 => "011010100100001010100",
		348 => "011010100100001110100",
		349 => "011010100100001110100",
		350 => "011010100100001110100",
		351 => "011000001101100010011",
		352 => "011000001101100010011",
		353 => "011000001101100010011",
		354 => "011000001101100010011",
		355 => "011000001101100010011",
		356 => "011000001101100010011",
		357 => "011010100100001010100",
		358 => "011010100100001010100",
		359 => "011010100100001010100",
		360 => "011010100100001110100",
		361 => "011010100100001110100",
		362 => "011010100100001110100",
		363 => "011000001101100010011",
		364 => "011000001101100010011",
		365 => "011000001101100010011",
		366 => "111011010100001010011",
		367 => "111011010100001010011",
		368 => "111011010100001010011",
		369 => "011010100100001010100",
		370 => "011010100100001010100",
		371 => "011010100100001010100",
		372 => "011010100100001110100",
		373 => "011010100100001110100",
		374 => "011010100100001110100",
		375 => "011000001101100010011",
		376 => "011000001101100010011",
		377 => "011000001101100010011",
		378 => "011000001101100010011",
		379 => "011000001101100010011",
		380 => "011000001101100010011",
		381 => "011010100100001010100",
		382 => "011010100100001010100",
		383 => "011010100100001010100",
		384 => "011001111100001010110",
		385 => "011001111100001010110",
		386 => "011001111100001010110",
		387 => "011001100100001110001",
		388 => "011001100100001110001",
		389 => "011001100100001110001",
		390 => "011011000100001110011",
		391 => "011011000100001110011",
		392 => "011011000100001110011",
		393 => "001000111100111010000",
		394 => "001000111100111010000",
		395 => "001000111100111010000",
		396 => "011001111100001010110",
		397 => "011001111100001010110",
		398 => "011001111100001010110",
		399 => "011001100100001110001",
		400 => "011001100100001110001",
		401 => "011001100100001110001",
		402 => "011011000100001110011",
		403 => "011011000100001110011",
		404 => "011011000100001110011",
		405 => "001000111100111010000",
		406 => "001000111100111010000",
		407 => "001000111100111010000",
		408 => "011001111100001010110",
		409 => "011001111100001010110",
		410 => "011001111100001010110",
		411 => "011001100100001110001",
		412 => "011001100100001110001",
		413 => "011001100100001110001",
		414 => "011011000100001110011",
		415 => "011011000100001110011",
		416 => "011011000100001110011",
		417 => "001000111100111010000",
		418 => "001000111100111010000",
		419 => "001000111100111010000",
		420 => "011001111100001010110",
		421 => "011001111100001010110",
		422 => "011001111100001010110",
		423 => "011001100100001110001",
		424 => "011001100100001110001",
		425 => "011001100100001110001",
		426 => "011011000100001110011",
		427 => "011011000100001110011",
		428 => "011011000100001110011",
		429 => "001000111100111010000",
		430 => "001000111100111010000",
		431 => "001000111100111010000",
		432 => "011001111100001010110",
		433 => "011001111100001010110",
		434 => "011001111100001010110",
		435 => "011001100100001110001",
		436 => "011001100100001110001",
		437 => "011001100100001110001",
		438 => "011011000100001110011",
		439 => "011011000100001110011",
		440 => "011011000100001110011",
		441 => "001000111100111010000",
		442 => "001000111100111010000",
		443 => "001000111100111010000",
		444 => "011001111100001010110",
		445 => "011001111100001010110",
		446 => "011001111100001010110",
		447 => "011001100100001110001",
		448 => "011001100100001110001",
		449 => "011001100100001110001",
		450 => "011011000100001110011",
		451 => "011011000100001110011",
		452 => "011011000100001110011",
		453 => "001000111100111010000",
		454 => "001000111100111010000",
		455 => "001000111100111010000",
		456 => "011001111100001010110",
		457 => "011001111100001010110",
		458 => "011001111100001010110",
		459 => "011001100100001110001",
		460 => "011001100100001110001",
		461 => "011001100100001110001",
		462 => "011011000100001110011",
		463 => "011011000100001110011",
		464 => "011011000100001110011",
		465 => "001000111100111010000",
		466 => "001000111100111010000",
		467 => "001000111100111010000",
		468 => "011001111100001010110",
		469 => "011001111100001010110",
		470 => "011001111100001010110",
		471 => "011001100100001110001",
		472 => "011001100100001110001",
		473 => "011001100100001110001",
		474 => "011011000100001110011",
		475 => "011011000100001110011",
		476 => "011011000100001110011",
		477 => "001000111100111010000",
		478 => "001000111100111010000",
		479 => "001000111100111010000",
		480 => "011000101100100010101",
		481 => "011000101100100010101",
		482 => "011000101100100010101",
		483 => "011000101100100010101",
		484 => "011000101100100010101",
		485 => "011000101100100010101",
		486 => "011000101100100010101",
		487 => "011000101100100010101",
		488 => "011000101100100010101",
		489 => "011000101100100010101",
		490 => "011000101100100010101",
		491 => "011000101100100010101",
		492 => "011000101100100010101",
		493 => "011000101100100010101",
		494 => "011000101100100010101",
		495 => "011000101100100010101",
		496 => "011000101100100010101",
		497 => "011000101100100010101",
		498 => "011000101100100010101",
		499 => "011000101100100010101",
		500 => "011000101100100010101",
		501 => "011000101100100010101",
		502 => "011000101100100010101",
		503 => "011000101100100010101",
		504 => "011000101100100010101",
		505 => "011000101100100010101",
		506 => "011000101100100010101",
		507 => "011000101100100010101",
		508 => "011000101100100010101",
		509 => "011000101100100010101",
		510 => "011000101100100010101",
		511 => "011000101100100010101",
		512 => "011000101100100010101",
		513 => "011000101100100010101",
		514 => "011000101100100010101",
		515 => "011000101100100010101",
		516 => "011000101100100010101",
		517 => "011000101100100010101",
		518 => "011000101100100010101",
		519 => "011000101100100010101",
		520 => "011000101100100010101",
		521 => "011000101100100010101",
		522 => "011000101100100010101",
		523 => "011000101100100010101",
		524 => "011000101100100010101",
		525 => "011000101100100010101",
		526 => "011000101100100010101",
		527 => "011000101100100010101",
		528 => "011000101100100010101",
		529 => "011000101100100010101",
		530 => "011000101100100010101",
		531 => "011000101100100010101",
		532 => "011000101100100010101",
		533 => "011000101100100010101",
		534 => "011000101100100010101",
		535 => "011000101100100010101",
		536 => "011000101100100010101",
		537 => "011000101100100010101",
		538 => "011000101100100010101",
		539 => "011000101100100010101",
		540 => "011000101100100010101",
		541 => "011000101100100010101",
		542 => "011000101100100010101",
		543 => "011000101100100010101",
		544 => "011000101100100010101",
		545 => "011000101100100010101",
		546 => "011000101100100010101",
		547 => "011000101100100010101",
		548 => "011000101100100010101",
		549 => "011000101100100010101",
		550 => "011000101100100010101",
		551 => "011000101100100010101",
		552 => "011000101100100010101",
		553 => "011000101100100010101",
		554 => "011000101100100010101",
		555 => "011000101100100010101",
		556 => "011000101100100010101",
		557 => "011000101100100010101",
		558 => "011000101100100010101",
		559 => "011000101100100010101",
		560 => "011000101100100010101",
		561 => "011000101100100010101",
		562 => "011000101100100010101",
		563 => "011000101100100010101",
		564 => "011000101100100010101",
		565 => "011000101100100010101",
		566 => "011000101100100010101",
		567 => "011000101100100010101",
		568 => "011000101100100010101",
		569 => "011000101100100010101",
		570 => "011000101100100010101",
		571 => "011000101100100010101",
		572 => "011000101100100010101",
		573 => "011000101100100010101",
		574 => "011000101100100010101",
		575 => "011000101100100010101",
		576 => "011000101100100110010",
		577 => "011000101100100110010",
		578 => "011000101100100110010",
		579 => "011000101100100110010",
		580 => "011000101100100110010",
		581 => "011000101100100110010",
		582 => "011000101100100110010",
		583 => "011000101100100110010",
		584 => "011000101100100110010",
		585 => "011000101100100110010",
		586 => "011000101100100110010",
		587 => "011000101100100110010",
		588 => "011000101100100110010",
		589 => "011000101100100110010",
		590 => "011000101100100110010",
		591 => "011000101100100110010",
		592 => "011000101100100110010",
		593 => "011000101100100110010",
		594 => "011000101100100110010",
		595 => "011000101100100110010",
		596 => "011000101100100110010",
		597 => "011000101100100110010",
		598 => "011000101100100110010",
		599 => "011000101100100110010",
		600 => "011000101100100110010",
		601 => "011000101100100110010",
		602 => "011000101100100110010",
		603 => "011000101100100110010",
		604 => "011000101100100110010",
		605 => "011000101100100110010",
		606 => "011000101100100110010",
		607 => "011000101100100110010",
		608 => "011000101100100110010",
		609 => "011000101100100110010",
		610 => "011000101100100110010",
		611 => "011000101100100110010",
		612 => "011000101100100110010",
		613 => "011000101100100110010",
		614 => "011000101100100110010",
		615 => "011000101100100110010",
		616 => "011000101100100110010",
		617 => "011000101100100110010",
		618 => "011000101100100110010",
		619 => "011000101100100110010",
		620 => "011000101100100110010",
		621 => "011000101100100110010",
		622 => "011000101100100110010",
		623 => "011000101100100110010",
		624 => "011000101100100110010",
		625 => "011000101100100110010",
		626 => "011000101100100110010",
		627 => "011000101100100110010",
		628 => "011000101100100110010",
		629 => "011000101100100110010",
		630 => "011000101100100110010",
		631 => "011000101100100110010",
		632 => "011000101100100110010",
		633 => "011000101100100110010",
		634 => "011000101100100110010",
		635 => "011000101100100110010",
		636 => "011000101100100110010",
		637 => "011000101100100110010",
		638 => "011000101100100110010",
		639 => "011000101100100110010",
		640 => "011000101100100110010",
		641 => "011000101100100110010",
		642 => "011000101100100110010",
		643 => "011000101100100110010",
		644 => "011000101100100110010",
		645 => "011000101100100110010",
		646 => "011000101100100110010",
		647 => "011000101100100110010",
		648 => "011000101100100110010",
		649 => "011000101100100110010",
		650 => "011000101100100110010",
		651 => "011000101100100110010",
		652 => "011000101100100110010",
		653 => "011000101100100110010",
		654 => "011000101100100110010",
		655 => "011000101100100110010",
		656 => "011000101100100110010",
		657 => "011000101100100110010",
		658 => "011000101100100110010",
		659 => "011000101100100110010",
		660 => "011000101100100110010",
		661 => "011000101100100110010",
		662 => "011000101100100110010",
		663 => "011000101100100110010",
		664 => "011000101100100110010",
		665 => "011000101100100110010",
		666 => "011000101100100110010",
		667 => "011000101100100110010",
		668 => "011000101100100110010",
		669 => "011000101100100110010",
		670 => "011000101100100110010",
		671 => "011000101100100110010",
		672 => "111000010100001010000",
		673 => "111000010100001010000",
		674 => "111000010100001010000",
		675 => "111000010100001010000",
		676 => "111000010100001010000",
		677 => "111000010100001010000",
		678 => "111000010100001010000",
		679 => "111000010100001010000",
		680 => "111000010100001010000",
		681 => "111000010100001010000",
		682 => "111000010100001010000",
		683 => "111000010100001010000",
		684 => "111000010100001010000",
		685 => "111000010100001010000",
		686 => "111000010100001010000",
		687 => "111000010100001010000",
		688 => "111000010100001010000",
		689 => "111000010100001010000",
		690 => "111000010100001010000",
		691 => "111000010100001010000",
		692 => "111000010100001010000",
		693 => "111000010100001010000",
		694 => "111000010100001010000",
		695 => "111000010100001010000",
		696 => "111000010100001010000",
		697 => "111000010100001010000",
		698 => "111000010100001010000",
		699 => "111000010100001010000",
		700 => "111000010100001010000",
		701 => "111000010100001010000",
		702 => "111000010100001010000",
		703 => "111000010100001010000",
		704 => "111000010100001010000",
		705 => "111000010100001010000",
		706 => "111000010100001010000",
		707 => "111000010100001010000",
		708 => "111000010100001010000",
		709 => "111000010100001010000",
		710 => "111000010100001010000",
		711 => "111000010100001010000",
		712 => "111000010100001010000",
		713 => "111000010100001010000",
		714 => "111000010100001010000",
		715 => "111000010100001010000",
		716 => "111000010100001010000",
		717 => "111000010100001010000",
		718 => "111000010100001010000",
		719 => "111000010100001010000",
		720 => "111000010100001010000",
		721 => "111000010100001010000",
		722 => "111000010100001010000",
		723 => "111000010100001010000",
		724 => "111000010100001010000",
		725 => "111000010100001010000",
		726 => "111000010100001010000",
		727 => "111000010100001010000",
		728 => "111000010100001010000",
		729 => "111000010100001010000",
		730 => "111000010100001010000",
		731 => "111000010100001010000",
		732 => "111000010100001010000",
		733 => "111000010100001010000",
		734 => "111000010100001010000",
		735 => "111000010100001010000",
		736 => "111000010100001010000",
		737 => "111000010100001010000",
		738 => "111000010100001010000",
		739 => "111000010100001010000",
		740 => "111000010100001010000",
		741 => "111000010100001010000",
		742 => "111000010100001010000",
		743 => "111000010100001010000",
		744 => "111000010100001010000",
		745 => "111000010100001010000",
		746 => "111000010100001010000",
		747 => "111000010100001010000",
		748 => "111000010100001010000",
		749 => "111000010100001010000",
		750 => "111000010100001010000",
		751 => "111000010100001010000",
		752 => "111000010100001010000",
		753 => "111000010100001010000",
		754 => "111000010100001010000",
		755 => "111000010100001010000",
		756 => "111000010100001010000",
		757 => "111000010100001010000",
		758 => "111000010100001010000",
		759 => "111000010100001010000",
		760 => "111000010100001010000",
		761 => "111000010100001010000",
		762 => "111000010100001010000",
		763 => "111000010100001010000",
		764 => "111000010100001010000",
		765 => "111000010100001010000",
		766 => "111000010100001010000",
		767 => "111000010100001010000",
		768 => "111000010100001010000",
		769 => "111000010100001010000",
		770 => "111000010100001010000",
		771 => "111000010100001010000",
		772 => "111000010100001010000",
		773 => "111000010100001010000",
		774 => "111000010100001010000",
		775 => "111000010100001010000",
		776 => "111000010100001010000",
		777 => "111000010100001010000",
		778 => "111000010100001010000",
		779 => "111000010100001010000",
		780 => "111000010100001010000",
		781 => "111000010100001010000",
		782 => "111000010100001010000",
		783 => "111000010100001010000",
		784 => "111000010100001010000",
		785 => "111000010100001010000",
		786 => "111000010100001010000",
		787 => "111000010100001010000",
		788 => "111000010100001010000",
		789 => "111000010100001010000",
		790 => "111000010100001010000",
		791 => "111000010100001010000",
		792 => "111000010100001010000",
		793 => "111000010100001010000",
		794 => "111000010100001010000",
		795 => "111000010100001010000",
		796 => "111000010100001010000",
		797 => "111000010100001010000",
		798 => "111000010100001010000",
		799 => "111000010100001010000",
		800 => "111000010100001010000",
		801 => "111000010100001010000",
		802 => "111000010100001010000",
		803 => "111000010100001010000",
		804 => "111000010100001010000",
		805 => "111000010100001010000",
		806 => "111000010100001010000",
		807 => "111000010100001010000",
		808 => "111000010100001010000",
		809 => "111000010100001010000",
		810 => "111000010100001010000",
		811 => "111000010100001010000",
		812 => "111000010100001010000",
		813 => "111000010100001010000",
		814 => "111000010100001010000",
		815 => "111000010100001010000",
		816 => "111000010100001010000",
		817 => "111000010100001010000",
		818 => "111000010100001010000",
		819 => "111000010100001010000",
		820 => "111000010100001010000",
		821 => "111000010100001010000",
		822 => "111000010100001010000",
		823 => "111000010100001010000",
		824 => "111000010100001010000",
		825 => "111000010100001010000",
		826 => "111000010100001010000",
		827 => "111000010100001010000",
		828 => "111000010100001010000",
		829 => "111000010100001010000",
		830 => "111000010100001010000",
		831 => "111000010100001010000",
		832 => "111000010100001010000",
		833 => "111000010100001010000",
		834 => "111000010100001010000",
		835 => "111000010100001010000",
		836 => "111000010100001010000",
		837 => "111000010100001010000",
		838 => "111000010100001010000",
		839 => "111000010100001010000",
		840 => "111000010100001010000",
		841 => "111000010100001010000",
		842 => "111000010100001010000",
		843 => "111000010100001010000",
		844 => "111000010100001010000",
		845 => "111000010100001010000",
		846 => "111000010100001010000",
		847 => "111000010100001010000",
		848 => "111000010100001010000",
		849 => "111000010100001010000",
		850 => "111000010100001010000",
		851 => "111000010100001010000",
		852 => "111000010100001010000",
		853 => "111000010100001010000",
		854 => "111000010100001010000",
		855 => "111000010100001010000",
		856 => "111000010100001010000",
		857 => "111000010100001010000",
		858 => "111000010100001010000",
		859 => "111000010100001010000",
		860 => "111000010100001010000",
		861 => "111000010100001010000",
		862 => "111000010100001010000",
		863 => "111000010100001010000");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;