library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT12 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT12;

architecture Behavioral of ROMFFT12 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 13 
	constant ROM_tb : ROM := (
		0 => "011011101110001010000",
		1 => "011011101110001010000",
		2 => "011011101110001010000",
		3 => "001010011100001010111",
		4 => "001010011100001010111",
		5 => "001010011100001010111",
		6 => "001001100101101110000",
		7 => "001001100101101110000",
		8 => "001001100101101110000",
		9 => "011010100100001010010",
		10 => "011010100100001010010",
		11 => "011010100100001010010",
		12 => "011000001101100010011",
		13 => "011000001101100010011",
		14 => "011000001101100010011",
		15 => "001001011100001010100",
		16 => "001001011100001010100",
		17 => "001001011100001010100",
		18 => "011000001100101010110",
		19 => "011000001100101010110",
		20 => "011000001100101010110",
		21 => "011000011100111010000",
		22 => "011000011100111010000",
		23 => "011000011100111010000",
		24 => "011000101100101010100",
		25 => "011000101100101010100",
		26 => "011000101100101010100",
		27 => "001001111100011110010",
		28 => "001001111100011110010",
		29 => "001001111100011110010",
		30 => "011000000100111010001",
		31 => "011000000100111010001",
		32 => "011000000100111010001",
		33 => "001000110100001010011",
		34 => "001000110100001010011",
		35 => "001000110100001010011",
		36 => "011000000101011010010",
		37 => "011000000101011010010",
		38 => "011000000101011010010",
		39 => "011000000101011010010",
		40 => "011000000101011010010",
		41 => "011000000101011010010",
		42 => "001001111110001010000",
		43 => "001001111110001010000",
		44 => "001001111110001010000",
		45 => "011000000110111010101",
		46 => "011000000110111010101",
		47 => "011000000110111010101",
		48 => "001000011110001010110",
		49 => "001000011110001010110",
		50 => "001000011110001010110",
		51 => "001000011101101010011",
		52 => "001000011101101010011",
		53 => "001000011101101010011",
		54 => "001000010100111010110",
		55 => "001000010100111010110",
		56 => "001000010100111010110",
		57 => "011010100100001010010",
		58 => "011010100100001010010",
		59 => "011010100100001010010",
		60 => "011000001101100010011",
		61 => "011000001101100010011",
		62 => "011000001101100010011",
		63 => "011010000100001010010",
		64 => "011010000100001010010",
		65 => "011010000100001010010",
		66 => "001000111100011110011",
		67 => "001000111100011110011",
		68 => "001000111100011110011",
		69 => "011001000100001110100",
		70 => "011001000100001110100",
		71 => "011001000100001110100",
		72 => "011001000100001110100",
		73 => "011001000100001110100",
		74 => "011001000100001110100",
		75 => "011001000100001010011",
		76 => "011001000100001010011",
		77 => "011001000100001010011",
		78 => "011000000100111010001",
		79 => "011000000100111010001",
		80 => "011000000100111010001",
		81 => "011000101100100110100",
		82 => "011000101100100110100",
		83 => "011000101100100110100",
		84 => "011000000101011010010",
		85 => "011000000101011010010",
		86 => "011000000101011010010",
		87 => "001001011101011010000",
		88 => "001001011101011010000",
		89 => "001001011101011010000",
		90 => "001001111110001010000",
		91 => "001001111110001010000",
		92 => "001001111110001010000",
		93 => "001000011110101010111",
		94 => "001000011110101010111",
		95 => "001000011110101010111",
		96 => "011000000101110011001",
		97 => "011000000101110011001",
		98 => "011000000101110011001",
		99 => "001001111100001010101",
		100 => "001001111100001010101",
		101 => "001001111100001010101",
		102 => "001011011100001010111",
		103 => "001011011100001010111",
		104 => "001011011100001010111",
		105 => "011001011100111010000",
		106 => "011001011100111010000",
		107 => "011001011100111010000",
		108 => "011000000101101010011",
		109 => "011000000101101010011",
		110 => "011000000101101010011",
		111 => "011000001101110010011",
		112 => "011000001101110010011",
		113 => "011000001101110010011",
		114 => "011000001110100010101",
		115 => "011000001110100010101",
		116 => "011000001110100010101",
		117 => "011000000110011010100",
		118 => "011000000110011010100",
		119 => "011000000110011010100",
		120 => "011000000101110011001",
		121 => "011000000101110011001",
		122 => "011000000101110011001",
		123 => "001000011101011010010",
		124 => "001000011101011010010",
		125 => "001000011101011010010",
		126 => "011000111100111010000",
		127 => "011000111100111010000",
		128 => "011000111100111010000",
		129 => "011001100100001010010",
		130 => "011001100100001010010",
		131 => "011001100100001010010",
		132 => "011000000101101010011",
		133 => "011000000101101010011",
		134 => "011000000101101010011",
		135 => "011000001101110010011",
		136 => "011000001101110010011",
		137 => "011000001101110010011",
		138 => "011000001110100010101",
		139 => "011000001110100010101",
		140 => "011000001110100010101",
		141 => "001010011110011010000",
		142 => "001010011110011010000",
		143 => "001010011110011010000",
		144 => "011000000101110011001",
		145 => "011000000101110011001",
		146 => "011000000101110011001",
		147 => "001001111100001010101",
		148 => "001001111100001010101",
		149 => "001001111100001010101",
		150 => "001011011100001010111",
		151 => "001011011100001010111",
		152 => "001011011100001010111",
		153 => "011001011100111010000",
		154 => "011001011100111010000",
		155 => "011001011100111010000",
		156 => "011000000101101010011",
		157 => "011000000101101010011",
		158 => "011000000101101010011",
		159 => "011000001101110010011",
		160 => "011000001101110010011",
		161 => "011000001101110010011",
		162 => "011000001110100010101",
		163 => "011000001110100010101",
		164 => "011000001110100010101",
		165 => "011000000110011010100",
		166 => "011000000110011010100",
		167 => "011000000110011010100",
		168 => "011000000101110011001",
		169 => "011000000101110011001",
		170 => "011000000101110011001",
		171 => "001000011101011010010",
		172 => "001000011101011010010",
		173 => "001000011101011010010",
		174 => "011000111100111010000",
		175 => "011000111100111010000",
		176 => "011000111100111010000",
		177 => "011001100100001010010",
		178 => "011001100100001010010",
		179 => "011001100100001010010",
		180 => "011000000101101010011",
		181 => "011000000101101010011",
		182 => "011000000101101010011",
		183 => "011000001101110010011",
		184 => "011000001101110010011",
		185 => "011000001101110010011",
		186 => "011000001110100010101",
		187 => "011000001110100010101",
		188 => "011000001110100010101",
		189 => "001010011110011010000",
		190 => "001010011110011010000",
		191 => "001010011110011010000",
		192 => "001010111100001010101",
		193 => "001010111100001010101",
		194 => "001010111100001010101",
		195 => "001000111100011110011",
		196 => "001000111100011110011",
		197 => "001000111100011110011",
		198 => "011001011100001010100",
		199 => "011001011100001010100",
		200 => "011001011100001010100",
		201 => "011011100100001110011",
		202 => "011011100100001110011",
		203 => "011011100100001110011",
		204 => "011010100100001010101",
		205 => "011010100100001010101",
		206 => "011010100100001010101",
		207 => "001000100100111010001",
		208 => "001000100100111010001",
		209 => "001000100100111010001",
		210 => "011010000100001110010",
		211 => "011010000100001110010",
		212 => "011010000100001110010",
		213 => "011000000101111010011",
		214 => "011000000101111010011",
		215 => "011000000101111010011",
		216 => "001010111100001010101",
		217 => "001010111100001010101",
		218 => "001010111100001010101",
		219 => "001000111100011110011",
		220 => "001000111100011110011",
		221 => "001000111100011110011",
		222 => "011001011100001010100",
		223 => "011001011100001010100",
		224 => "011001011100001010100",
		225 => "011011100100001110011",
		226 => "011011100100001110011",
		227 => "011011100100001110011",
		228 => "011010100100001010101",
		229 => "011010100100001010101",
		230 => "011010100100001010101",
		231 => "001000100100111010001",
		232 => "001000100100111010001",
		233 => "001000100100111010001",
		234 => "011010000100001110010",
		235 => "011010000100001110010",
		236 => "011010000100001110010",
		237 => "011000000101111010011",
		238 => "011000000101111010011",
		239 => "011000000101111010011",
		240 => "001010111100001010101",
		241 => "001010111100001010101",
		242 => "001010111100001010101",
		243 => "001000111100011110011",
		244 => "001000111100011110011",
		245 => "001000111100011110011",
		246 => "011001011100001010100",
		247 => "011001011100001010100",
		248 => "011001011100001010100",
		249 => "011011100100001110011",
		250 => "011011100100001110011",
		251 => "011011100100001110011",
		252 => "011010100100001010101",
		253 => "011010100100001010101",
		254 => "011010100100001010101",
		255 => "001000100100111010001",
		256 => "001000100100111010001",
		257 => "001000100100111010001",
		258 => "011010000100001110010",
		259 => "011010000100001110010",
		260 => "011010000100001110010",
		261 => "011000000101111010011",
		262 => "011000000101111010011",
		263 => "011000000101111010011",
		264 => "001010111100001010101",
		265 => "001010111100001010101",
		266 => "001010111100001010101",
		267 => "001000111100011110011",
		268 => "001000111100011110011",
		269 => "001000111100011110011",
		270 => "011001011100001010100",
		271 => "011001011100001010100",
		272 => "011001011100001010100",
		273 => "011011100100001110011",
		274 => "011011100100001110011",
		275 => "011011100100001110011",
		276 => "011010100100001010101",
		277 => "011010100100001010101",
		278 => "011010100100001010101",
		279 => "001000100100111010001",
		280 => "001000100100111010001",
		281 => "001000100100111010001",
		282 => "011010000100001110010",
		283 => "011010000100001110010",
		284 => "011010000100001110010",
		285 => "011000000101111010011",
		286 => "011000000101111010011",
		287 => "011000000101111010011",
		288 => "011000001101100010011",
		289 => "011000001101100010011",
		290 => "011000001101100010011",
		291 => "011010100100001010100",
		292 => "011010100100001010100",
		293 => "011010100100001010100",
		294 => "011000001101100010011",
		295 => "011000001101100010011",
		296 => "011000001101100010011",
		297 => "011010100100001010100",
		298 => "011010100100001010100",
		299 => "011010100100001010100",
		300 => "011000001101100010011",
		301 => "011000001101100010011",
		302 => "011000001101100010011",
		303 => "011010100100001010100",
		304 => "011010100100001010100",
		305 => "011010100100001010100",
		306 => "011000001101100010011",
		307 => "011000001101100010011",
		308 => "011000001101100010011",
		309 => "011010100100001010100",
		310 => "011010100100001010100",
		311 => "011010100100001010100",
		312 => "011000001101100010011",
		313 => "011000001101100010011",
		314 => "011000001101100010011",
		315 => "011010100100001010100",
		316 => "011010100100001010100",
		317 => "011010100100001010100",
		318 => "011000001101100010011",
		319 => "011000001101100010011",
		320 => "011000001101100010011",
		321 => "011010100100001010100",
		322 => "011010100100001010100",
		323 => "011010100100001010100",
		324 => "011000001101100010011",
		325 => "011000001101100010011",
		326 => "011000001101100010011",
		327 => "011010100100001010100",
		328 => "011010100100001010100",
		329 => "011010100100001010100",
		330 => "011000001101100010011",
		331 => "011000001101100010011",
		332 => "011000001101100010011",
		333 => "011010100100001010100",
		334 => "011010100100001010100",
		335 => "011010100100001010100",
		336 => "011000001101100010011",
		337 => "011000001101100010011",
		338 => "011000001101100010011",
		339 => "011010100100001010100",
		340 => "011010100100001010100",
		341 => "011010100100001010100",
		342 => "011000001101100010011",
		343 => "011000001101100010011",
		344 => "011000001101100010011",
		345 => "011010100100001010100",
		346 => "011010100100001010100",
		347 => "011010100100001010100",
		348 => "011000001101100010011",
		349 => "011000001101100010011",
		350 => "011000001101100010011",
		351 => "011010100100001010100",
		352 => "011010100100001010100",
		353 => "011010100100001010100",
		354 => "011000001101100010011",
		355 => "011000001101100010011",
		356 => "011000001101100010011",
		357 => "011010100100001010100",
		358 => "011010100100001010100",
		359 => "011010100100001010100",
		360 => "011000001101100010011",
		361 => "011000001101100010011",
		362 => "011000001101100010011",
		363 => "011010100100001010100",
		364 => "011010100100001010100",
		365 => "011010100100001010100",
		366 => "011000001101100010011",
		367 => "011000001101100010011",
		368 => "011000001101100010011",
		369 => "011010100100001010100",
		370 => "011010100100001010100",
		371 => "011010100100001010100",
		372 => "011000001101100010011",
		373 => "011000001101100010011",
		374 => "011000001101100010011",
		375 => "011010100100001010100",
		376 => "011010100100001010100",
		377 => "011010100100001010100",
		378 => "011000001101100010011",
		379 => "011000001101100010011",
		380 => "011000001101100010011",
		381 => "011010100100001010100",
		382 => "011010100100001010100",
		383 => "011010100100001010100",
		384 => "011001100100001110001",
		385 => "011001100100001110001",
		386 => "011001100100001110001",
		387 => "001000111100111010000",
		388 => "001000111100111010000",
		389 => "001000111100111010000",
		390 => "011001100100001110001",
		391 => "011001100100001110001",
		392 => "011001100100001110001",
		393 => "001000111100111010000",
		394 => "001000111100111010000",
		395 => "001000111100111010000",
		396 => "011001100100001110001",
		397 => "011001100100001110001",
		398 => "011001100100001110001",
		399 => "001000111100111010000",
		400 => "001000111100111010000",
		401 => "001000111100111010000",
		402 => "011001100100001110001",
		403 => "011001100100001110001",
		404 => "011001100100001110001",
		405 => "001000111100111010000",
		406 => "001000111100111010000",
		407 => "001000111100111010000",
		408 => "011001100100001110001",
		409 => "011001100100001110001",
		410 => "011001100100001110001",
		411 => "001000111100111010000",
		412 => "001000111100111010000",
		413 => "001000111100111010000",
		414 => "011001100100001110001",
		415 => "011001100100001110001",
		416 => "011001100100001110001",
		417 => "001000111100111010000",
		418 => "001000111100111010000",
		419 => "001000111100111010000",
		420 => "011001100100001110001",
		421 => "011001100100001110001",
		422 => "011001100100001110001",
		423 => "001000111100111010000",
		424 => "001000111100111010000",
		425 => "001000111100111010000",
		426 => "011001100100001110001",
		427 => "011001100100001110001",
		428 => "011001100100001110001",
		429 => "001000111100111010000",
		430 => "001000111100111010000",
		431 => "001000111100111010000",
		432 => "011001100100001110001",
		433 => "011001100100001110001",
		434 => "011001100100001110001",
		435 => "001000111100111010000",
		436 => "001000111100111010000",
		437 => "001000111100111010000",
		438 => "011001100100001110001",
		439 => "011001100100001110001",
		440 => "011001100100001110001",
		441 => "001000111100111010000",
		442 => "001000111100111010000",
		443 => "001000111100111010000",
		444 => "011001100100001110001",
		445 => "011001100100001110001",
		446 => "011001100100001110001",
		447 => "001000111100111010000",
		448 => "001000111100111010000",
		449 => "001000111100111010000",
		450 => "011001100100001110001",
		451 => "011001100100001110001",
		452 => "011001100100001110001",
		453 => "001000111100111010000",
		454 => "001000111100111010000",
		455 => "001000111100111010000",
		456 => "011001100100001110001",
		457 => "011001100100001110001",
		458 => "011001100100001110001",
		459 => "001000111100111010000",
		460 => "001000111100111010000",
		461 => "001000111100111010000",
		462 => "011001100100001110001",
		463 => "011001100100001110001",
		464 => "011001100100001110001",
		465 => "001000111100111010000",
		466 => "001000111100111010000",
		467 => "001000111100111010000",
		468 => "011001100100001110001",
		469 => "011001100100001110001",
		470 => "011001100100001110001",
		471 => "001000111100111010000",
		472 => "001000111100111010000",
		473 => "001000111100111010000",
		474 => "011001100100001110001",
		475 => "011001100100001110001",
		476 => "011001100100001110001",
		477 => "001000111100111010000",
		478 => "001000111100111010000",
		479 => "001000111100111010000",
		480 => "011000101100100010101",
		481 => "011000101100100010101",
		482 => "011000101100100010101",
		483 => "011000101100100010101",
		484 => "011000101100100010101",
		485 => "011000101100100010101",
		486 => "011000101100100010101",
		487 => "011000101100100010101",
		488 => "011000101100100010101",
		489 => "011000101100100010101",
		490 => "011000101100100010101",
		491 => "011000101100100010101",
		492 => "011000101100100010101",
		493 => "011000101100100010101",
		494 => "011000101100100010101",
		495 => "011000101100100010101",
		496 => "011000101100100010101",
		497 => "011000101100100010101",
		498 => "011000101100100010101",
		499 => "011000101100100010101",
		500 => "011000101100100010101",
		501 => "011000101100100010101",
		502 => "011000101100100010101",
		503 => "011000101100100010101",
		504 => "011000101100100010101",
		505 => "011000101100100010101",
		506 => "011000101100100010101",
		507 => "011000101100100010101",
		508 => "011000101100100010101",
		509 => "011000101100100010101",
		510 => "011000101100100010101",
		511 => "011000101100100010101",
		512 => "011000101100100010101",
		513 => "011000101100100010101",
		514 => "011000101100100010101",
		515 => "011000101100100010101",
		516 => "011000101100100010101",
		517 => "011000101100100010101",
		518 => "011000101100100010101",
		519 => "011000101100100010101",
		520 => "011000101100100010101",
		521 => "011000101100100010101",
		522 => "011000101100100010101",
		523 => "011000101100100010101",
		524 => "011000101100100010101",
		525 => "011000101100100010101",
		526 => "011000101100100010101",
		527 => "011000101100100010101",
		528 => "011000101100100010101",
		529 => "011000101100100010101",
		530 => "011000101100100010101",
		531 => "011000101100100010101",
		532 => "011000101100100010101",
		533 => "011000101100100010101",
		534 => "011000101100100010101",
		535 => "011000101100100010101",
		536 => "011000101100100010101",
		537 => "011000101100100010101",
		538 => "011000101100100010101",
		539 => "011000101100100010101",
		540 => "011000101100100010101",
		541 => "011000101100100010101",
		542 => "011000101100100010101",
		543 => "011000101100100010101",
		544 => "011000101100100010101",
		545 => "011000101100100010101",
		546 => "011000101100100010101",
		547 => "011000101100100010101",
		548 => "011000101100100010101",
		549 => "011000101100100010101",
		550 => "011000101100100010101",
		551 => "011000101100100010101",
		552 => "011000101100100010101",
		553 => "011000101100100010101",
		554 => "011000101100100010101",
		555 => "011000101100100010101",
		556 => "011000101100100010101",
		557 => "011000101100100010101",
		558 => "011000101100100010101",
		559 => "011000101100100010101",
		560 => "011000101100100010101",
		561 => "011000101100100010101",
		562 => "011000101100100010101",
		563 => "011000101100100010101",
		564 => "011000101100100010101",
		565 => "011000101100100010101",
		566 => "011000101100100010101",
		567 => "011000101100100010101",
		568 => "011000101100100010101",
		569 => "011000101100100010101",
		570 => "011000101100100010101",
		571 => "011000101100100010101",
		572 => "011000101100100010101",
		573 => "011000101100100010101",
		574 => "011000101100100010101",
		575 => "011000101100100010101",
		576 => "011000101100100110010",
		577 => "011000101100100110010",
		578 => "011000101100100110010",
		579 => "011000101100100110010",
		580 => "011000101100100110010",
		581 => "011000101100100110010",
		582 => "011000101100100110010",
		583 => "011000101100100110010",
		584 => "011000101100100110010",
		585 => "011000101100100110010",
		586 => "011000101100100110010",
		587 => "011000101100100110010",
		588 => "011000101100100110010",
		589 => "011000101100100110010",
		590 => "011000101100100110010",
		591 => "011000101100100110010",
		592 => "011000101100100110010",
		593 => "011000101100100110010",
		594 => "011000101100100110010",
		595 => "011000101100100110010",
		596 => "011000101100100110010",
		597 => "011000101100100110010",
		598 => "011000101100100110010",
		599 => "011000101100100110010",
		600 => "011000101100100110010",
		601 => "011000101100100110010",
		602 => "011000101100100110010",
		603 => "011000101100100110010",
		604 => "011000101100100110010",
		605 => "011000101100100110010",
		606 => "011000101100100110010",
		607 => "011000101100100110010",
		608 => "011000101100100110010",
		609 => "011000101100100110010",
		610 => "011000101100100110010",
		611 => "011000101100100110010",
		612 => "011000101100100110010",
		613 => "011000101100100110010",
		614 => "011000101100100110010",
		615 => "011000101100100110010",
		616 => "011000101100100110010",
		617 => "011000101100100110010",
		618 => "011000101100100110010",
		619 => "011000101100100110010",
		620 => "011000101100100110010",
		621 => "011000101100100110010",
		622 => "011000101100100110010",
		623 => "011000101100100110010",
		624 => "011000101100100110010",
		625 => "011000101100100110010",
		626 => "011000101100100110010",
		627 => "011000101100100110010",
		628 => "011000101100100110010",
		629 => "011000101100100110010",
		630 => "011000101100100110010",
		631 => "011000101100100110010",
		632 => "011000101100100110010",
		633 => "011000101100100110010",
		634 => "011000101100100110010",
		635 => "011000101100100110010",
		636 => "011000101100100110010",
		637 => "011000101100100110010",
		638 => "011000101100100110010",
		639 => "011000101100100110010",
		640 => "011000101100100110010",
		641 => "011000101100100110010",
		642 => "011000101100100110010",
		643 => "011000101100100110010",
		644 => "011000101100100110010",
		645 => "011000101100100110010",
		646 => "011000101100100110010",
		647 => "011000101100100110010",
		648 => "011000101100100110010",
		649 => "011000101100100110010",
		650 => "011000101100100110010",
		651 => "011000101100100110010",
		652 => "011000101100100110010",
		653 => "011000101100100110010",
		654 => "011000101100100110010",
		655 => "011000101100100110010",
		656 => "011000101100100110010",
		657 => "011000101100100110010",
		658 => "011000101100100110010",
		659 => "011000101100100110010",
		660 => "011000101100100110010",
		661 => "011000101100100110010",
		662 => "011000101100100110010",
		663 => "011000101100100110010",
		664 => "011000101100100110010",
		665 => "011000101100100110010",
		666 => "011000101100100110010",
		667 => "011000101100100110010",
		668 => "011000101100100110010",
		669 => "011000101100100110010",
		670 => "011000101100100110010",
		671 => "011000101100100110010",
		672 => "111000010100001010000",
		673 => "111000010100001010000",
		674 => "111000010100001010000",
		675 => "111000010100001010000",
		676 => "111000010100001010000",
		677 => "111000010100001010000",
		678 => "111000010100001010000",
		679 => "111000010100001010000",
		680 => "111000010100001010000",
		681 => "111000010100001010000",
		682 => "111000010100001010000",
		683 => "111000010100001010000",
		684 => "111000010100001010000",
		685 => "111000010100001010000",
		686 => "111000010100001010000",
		687 => "111000010100001010000",
		688 => "111000010100001010000",
		689 => "111000010100001010000",
		690 => "111000010100001010000",
		691 => "111000010100001010000",
		692 => "111000010100001010000",
		693 => "111000010100001010000",
		694 => "111000010100001010000",
		695 => "111000010100001010000",
		696 => "111000010100001010000",
		697 => "111000010100001010000",
		698 => "111000010100001010000",
		699 => "111000010100001010000",
		700 => "111000010100001010000",
		701 => "111000010100001010000",
		702 => "111000010100001010000",
		703 => "111000010100001010000",
		704 => "111000010100001010000",
		705 => "111000010100001010000",
		706 => "111000010100001010000",
		707 => "111000010100001010000",
		708 => "111000010100001010000",
		709 => "111000010100001010000",
		710 => "111000010100001010000",
		711 => "111000010100001010000",
		712 => "111000010100001010000",
		713 => "111000010100001010000",
		714 => "111000010100001010000",
		715 => "111000010100001010000",
		716 => "111000010100001010000",
		717 => "111000010100001010000",
		718 => "111000010100001010000",
		719 => "111000010100001010000",
		720 => "111000010100001010000",
		721 => "111000010100001010000",
		722 => "111000010100001010000",
		723 => "111000010100001010000",
		724 => "111000010100001010000",
		725 => "111000010100001010000",
		726 => "111000010100001010000",
		727 => "111000010100001010000",
		728 => "111000010100001010000",
		729 => "111000010100001010000",
		730 => "111000010100001010000",
		731 => "111000010100001010000",
		732 => "111000010100001010000",
		733 => "111000010100001010000",
		734 => "111000010100001010000",
		735 => "111000010100001010000",
		736 => "111000010100001010000",
		737 => "111000010100001010000",
		738 => "111000010100001010000",
		739 => "111000010100001010000",
		740 => "111000010100001010000",
		741 => "111000010100001010000",
		742 => "111000010100001010000",
		743 => "111000010100001010000",
		744 => "111000010100001010000",
		745 => "111000010100001010000",
		746 => "111000010100001010000",
		747 => "111000010100001010000",
		748 => "111000010100001010000",
		749 => "111000010100001010000",
		750 => "111000010100001010000",
		751 => "111000010100001010000",
		752 => "111000010100001010000",
		753 => "111000010100001010000",
		754 => "111000010100001010000",
		755 => "111000010100001010000",
		756 => "111000010100001010000",
		757 => "111000010100001010000",
		758 => "111000010100001010000",
		759 => "111000010100001010000",
		760 => "111000010100001010000",
		761 => "111000010100001010000",
		762 => "111000010100001010000",
		763 => "111000010100001010000",
		764 => "111000010100001010000",
		765 => "111000010100001010000",
		766 => "111000010100001010000",
		767 => "111000010100001010000",
		768 => "111000010100001010000",
		769 => "111000010100001010000",
		770 => "111000010100001010000",
		771 => "111000010100001010000",
		772 => "111000010100001010000",
		773 => "111000010100001010000",
		774 => "111000010100001010000",
		775 => "111000010100001010000",
		776 => "111000010100001010000",
		777 => "111000010100001010000",
		778 => "111000010100001010000",
		779 => "111000010100001010000",
		780 => "111000010100001010000",
		781 => "111000010100001010000",
		782 => "111000010100001010000",
		783 => "111000010100001010000",
		784 => "111000010100001010000",
		785 => "111000010100001010000",
		786 => "111000010100001010000",
		787 => "111000010100001010000",
		788 => "111000010100001010000",
		789 => "111000010100001010000",
		790 => "111000010100001010000",
		791 => "111000010100001010000",
		792 => "111000010100001010000",
		793 => "111000010100001010000",
		794 => "111000010100001010000",
		795 => "111000010100001010000",
		796 => "111000010100001010000",
		797 => "111000010100001010000",
		798 => "111000010100001010000",
		799 => "111000010100001010000",
		800 => "111000010100001010000",
		801 => "111000010100001010000",
		802 => "111000010100001010000",
		803 => "111000010100001010000",
		804 => "111000010100001010000",
		805 => "111000010100001010000",
		806 => "111000010100001010000",
		807 => "111000010100001010000",
		808 => "111000010100001010000",
		809 => "111000010100001010000",
		810 => "111000010100001010000",
		811 => "111000010100001010000",
		812 => "111000010100001010000",
		813 => "111000010100001010000",
		814 => "111000010100001010000",
		815 => "111000010100001010000",
		816 => "111000010100001010000",
		817 => "111000010100001010000",
		818 => "111000010100001010000",
		819 => "111000010100001010000",
		820 => "111000010100001010000",
		821 => "111000010100001010000",
		822 => "111000010100001010000",
		823 => "111000010100001010000",
		824 => "111000010100001010000",
		825 => "111000010100001010000",
		826 => "111000010100001010000",
		827 => "111000010100001010000",
		828 => "111000010100001010000",
		829 => "111000010100001010000",
		830 => "111000010100001010000",
		831 => "111000010100001010000",
		832 => "111000010100001010000",
		833 => "111000010100001010000",
		834 => "111000010100001010000",
		835 => "111000010100001010000",
		836 => "111000010100001010000",
		837 => "111000010100001010000",
		838 => "111000010100001010000",
		839 => "111000010100001010000",
		840 => "111000010100001010000",
		841 => "111000010100001010000",
		842 => "111000010100001010000",
		843 => "111000010100001010000",
		844 => "111000010100001010000",
		845 => "111000010100001010000",
		846 => "111000010100001010000",
		847 => "111000010100001010000",
		848 => "111000010100001010000",
		849 => "111000010100001010000",
		850 => "111000010100001010000",
		851 => "111000010100001010000",
		852 => "111000010100001010000",
		853 => "111000010100001010000",
		854 => "111000010100001010000",
		855 => "111000010100001010000",
		856 => "111000010100001010000",
		857 => "111000010100001010000",
		858 => "111000010100001010000",
		859 => "111000010100001010000",
		860 => "111000010100001010000",
		861 => "111000010100001010000",
		862 => "111000010100001010000",
		863 => "111000010100001010000");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;