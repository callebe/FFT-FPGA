library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT10 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT10;

architecture Behavioral of ROMFFT10 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 11 
	constant ROM_tb : ROM := (
		0 => "001000011110101010100",
		1 => "001000011110101010100",
		2 => "001000011110101010100",
		3 => "011001111101111010000",
		4 => "011001111101111010000",
		5 => "011001111101111010000",
		6 => "001000010100101011000",
		7 => "001000010100101011000",
		8 => "001000010100101011000",
		9 => "011001001100111010000",
		10 => "011001001100111010000",
		11 => "011001001100111010000",
		12 => "011000001101010010011",
		13 => "011000001101010010011",
		14 => "011000001101010010011",
		15 => "011000111101001010000",
		16 => "011000111101001010000",
		17 => "011000111101001010000",
		18 => "001001111100001010110",
		19 => "001001111100001010110",
		20 => "001001111100001010110",
		21 => "001001011100001010011",
		22 => "001001011100001010011",
		23 => "001001011100001010011",
		24 => "011000000100111110000",
		25 => "011000000100111110000",
		26 => "011000000100111110000",
		27 => "001010011100011110010",
		28 => "001010011100011110010",
		29 => "001010011100011110010",
		30 => "011001100100001110001",
		31 => "011001100100001110001",
		32 => "011001100100001110001",
		33 => "011000000101001010100",
		34 => "011000000101001010100",
		35 => "011000000101001010100",
		36 => "011001100100001110001",
		37 => "011001100100001110001",
		38 => "011001100100001110001",
		39 => "011000000101101010010",
		40 => "011000000101101010010",
		41 => "011000000101101010010",
		42 => "011000000101111010011",
		43 => "011000000101111010011",
		44 => "011000000101111010011",
		45 => "011100001110011110000",
		46 => "011100001110011110000",
		47 => "011100001110011110000",
		48 => "011000001100110110110",
		49 => "011000001100110110110",
		50 => "011000001100110110110",
		51 => "011011100100001010011",
		52 => "011011100100001010011",
		53 => "011011100100001010011",
		54 => "011010100100001010111",
		55 => "011010100100001010111",
		56 => "011010100100001010111",
		57 => "011001100100011110000",
		58 => "011001100100011110000",
		59 => "011001100100011110000",
		60 => "011000001101010010011",
		61 => "011000001101010010011",
		62 => "011000001101010010011",
		63 => "011000111101001010000",
		64 => "011000111101001010000",
		65 => "011000111101001010000",
		66 => "011011000100001010011",
		67 => "011011000100001010011",
		68 => "011011000100001010011",
		69 => "011001100100001010010",
		70 => "011001100100001010010",
		71 => "011001100100001010010",
		72 => "001000011100001010011",
		73 => "001000011100001010011",
		74 => "001000011100001010011",
		75 => "011001000100001010100",
		76 => "011001000100001010100",
		77 => "011001000100001010100",
		78 => "001000111100111010000",
		79 => "001000111100111010000",
		80 => "001000111100111010000",
		81 => "011010000100001110100",
		82 => "011010000100001110100",
		83 => "011010000100001110100",
		84 => "001000111100111010000",
		85 => "001000111100111010000",
		86 => "001000111100111010000",
		87 => "011000000101101010010",
		88 => "011000000101101010010",
		89 => "011000000101101010010",
		90 => "011011100100001110011",
		91 => "011011100100001110011",
		92 => "011011100100001110011",
		93 => "001000011110001111001",
		94 => "001000011110001111001",
		95 => "001000011110001111001",
		96 => "011100000100001010011",
		97 => "011100000100001010011",
		98 => "011100000100001010011",
		99 => "001001011100001010101",
		100 => "001001011100001010101",
		101 => "001001011100001010101",
		102 => "011000000101111011000",
		103 => "011000000101111011000",
		104 => "011000000101111011000",
		105 => "001010011100011110010",
		106 => "001010011100011110010",
		107 => "001010011100011110010",
		108 => "001011011100001110010",
		109 => "001011011100001110010",
		110 => "001011011100001110010",
		111 => "011000001101100010011",
		112 => "011000001101100010011",
		113 => "011000001101100010011",
		114 => "011000000101101010011",
		115 => "011000000101101010011",
		116 => "011000000101101010011",
		117 => "011000011110001010110",
		118 => "011000011110001010110",
		119 => "011000011110001010110",
		120 => "011100000100001111001",
		121 => "011100000100001111001",
		122 => "011100000100001111001",
		123 => "011010100100001010010",
		124 => "011010100100001010010",
		125 => "011010100100001010010",
		126 => "001000111100001010011",
		127 => "001000111100001010011",
		128 => "001000111100001010011",
		129 => "011001000100001010100",
		130 => "011001000100001010100",
		131 => "011001000100001010100",
		132 => "001000000100101010110",
		133 => "001000000100101010110",
		134 => "001000000100101010110",
		135 => "011000001101100010011",
		136 => "011000001101100010011",
		137 => "011000001101100010011",
		138 => "001001100101101010000",
		139 => "001001100101101010000",
		140 => "001001100101101010000",
		141 => "011100000101101010000",
		142 => "011100000101101010000",
		143 => "011100000101101010000",
		144 => "011100000100001010011",
		145 => "011100000100001010011",
		146 => "011100000100001010011",
		147 => "001001011100001010101",
		148 => "001001011100001010101",
		149 => "001001011100001010101",
		150 => "011000000101111011000",
		151 => "011000000101111011000",
		152 => "011000000101111011000",
		153 => "001010011100011110010",
		154 => "001010011100011110010",
		155 => "001010011100011110010",
		156 => "001011011100001110010",
		157 => "001011011100001110010",
		158 => "001011011100001110010",
		159 => "011000001101100010011",
		160 => "011000001101100010011",
		161 => "011000001101100010011",
		162 => "011000000101101010011",
		163 => "011000000101101010011",
		164 => "011000000101101010011",
		165 => "011000011110001010110",
		166 => "011000011110001010110",
		167 => "011000011110001010110",
		168 => "011100000100001111001",
		169 => "011100000100001111001",
		170 => "011100000100001111001",
		171 => "011010100100001010010",
		172 => "011010100100001010010",
		173 => "011010100100001010010",
		174 => "001000111100001010011",
		175 => "001000111100001010011",
		176 => "001000111100001010011",
		177 => "011001000100001010100",
		178 => "011001000100001010100",
		179 => "011001000100001010100",
		180 => "001000000100101010110",
		181 => "001000000100101010110",
		182 => "001000000100101010110",
		183 => "011000001101100010011",
		184 => "011000001101100010011",
		185 => "011000001101100010011",
		186 => "001001100101101010000",
		187 => "001001100101101010000",
		188 => "001001100101101010000",
		189 => "011100000101101010000",
		190 => "011100000101101010000",
		191 => "011100000101101010000",
		192 => "011000001110100010101",
		193 => "011000001110100010101",
		194 => "011000001110100010101",
		195 => "001001111100001010110",
		196 => "001001111100001010110",
		197 => "001001111100001010110",
		198 => "011000111100001010011",
		199 => "011000111100001010011",
		200 => "011000111100001010011",
		201 => "011000010100111010110",
		202 => "011000010100111010110",
		203 => "011000010100111010110",
		204 => "011000001110100010101",
		205 => "011000001110100010101",
		206 => "011000001110100010101",
		207 => "011011000100001010011",
		208 => "011011000100001010011",
		209 => "011011000100001010011",
		210 => "011001100100001110001",
		211 => "011001100100001110001",
		212 => "011001100100001110001",
		213 => "011000000101110011001",
		214 => "011000000101110011001",
		215 => "011000000101110011001",
		216 => "011000001110100010101",
		217 => "011000001110100010101",
		218 => "011000001110100010101",
		219 => "001001111100001010110",
		220 => "001001111100001010110",
		221 => "001001111100001010110",
		222 => "011000111100001010011",
		223 => "011000111100001010011",
		224 => "011000111100001010011",
		225 => "011000010100111010110",
		226 => "011000010100111010110",
		227 => "011000010100111010110",
		228 => "011000001110100010101",
		229 => "011000001110100010101",
		230 => "011000001110100010101",
		231 => "011011000100001010011",
		232 => "011011000100001010011",
		233 => "011011000100001010011",
		234 => "011001100100001110001",
		235 => "011001100100001110001",
		236 => "011001100100001110001",
		237 => "011000000101110011001",
		238 => "011000000101110011001",
		239 => "011000000101110011001",
		240 => "011000001110100010101",
		241 => "011000001110100010101",
		242 => "011000001110100010101",
		243 => "001001111100001010110",
		244 => "001001111100001010110",
		245 => "001001111100001010110",
		246 => "011000111100001010011",
		247 => "011000111100001010011",
		248 => "011000111100001010011",
		249 => "011000010100111010110",
		250 => "011000010100111010110",
		251 => "011000010100111010110",
		252 => "011000001110100010101",
		253 => "011000001110100010101",
		254 => "011000001110100010101",
		255 => "011011000100001010011",
		256 => "011011000100001010011",
		257 => "011011000100001010011",
		258 => "011001100100001110001",
		259 => "011001100100001110001",
		260 => "011001100100001110001",
		261 => "011000000101110011001",
		262 => "011000000101110011001",
		263 => "011000000101110011001",
		264 => "011000001110100010101",
		265 => "011000001110100010101",
		266 => "011000001110100010101",
		267 => "001001111100001010110",
		268 => "001001111100001010110",
		269 => "001001111100001010110",
		270 => "011000111100001010011",
		271 => "011000111100001010011",
		272 => "011000111100001010011",
		273 => "011000010100111010110",
		274 => "011000010100111010110",
		275 => "011000010100111010110",
		276 => "011000001110100010101",
		277 => "011000001110100010101",
		278 => "011000001110100010101",
		279 => "011011000100001010011",
		280 => "011011000100001010011",
		281 => "011011000100001010011",
		282 => "011001100100001110001",
		283 => "011001100100001110001",
		284 => "011001100100001110001",
		285 => "011000000101110011001",
		286 => "011000000101110011001",
		287 => "011000000101110011001",
		288 => "011001011101001010000",
		289 => "011001011101001010000",
		290 => "011001011101001010000",
		291 => "011000000101011010101",
		292 => "011000000101011010101",
		293 => "011000000101011010101",
		294 => "011010000100001010010",
		295 => "011010000100001010010",
		296 => "011010000100001010010",
		297 => "011000000101011010101",
		298 => "011000000101011010101",
		299 => "011000000101011010101",
		300 => "011001011101001010000",
		301 => "011001011101001010000",
		302 => "011001011101001010000",
		303 => "011000000101011010101",
		304 => "011000000101011010101",
		305 => "011000000101011010101",
		306 => "011010000100001010010",
		307 => "011010000100001010010",
		308 => "011010000100001010010",
		309 => "011000000101011010101",
		310 => "011000000101011010101",
		311 => "011000000101011010101",
		312 => "011001011101001010000",
		313 => "011001011101001010000",
		314 => "011001011101001010000",
		315 => "011000000101011010101",
		316 => "011000000101011010101",
		317 => "011000000101011010101",
		318 => "011010000100001010010",
		319 => "011010000100001010010",
		320 => "011010000100001010010",
		321 => "011000000101011010101",
		322 => "011000000101011010101",
		323 => "011000000101011010101",
		324 => "011001011101001010000",
		325 => "011001011101001010000",
		326 => "011001011101001010000",
		327 => "011000000101011010101",
		328 => "011000000101011010101",
		329 => "011000000101011010101",
		330 => "011010000100001010010",
		331 => "011010000100001010010",
		332 => "011010000100001010010",
		333 => "011000000101011010101",
		334 => "011000000101011010101",
		335 => "011000000101011010101",
		336 => "011001011101001010000",
		337 => "011001011101001010000",
		338 => "011001011101001010000",
		339 => "011000000101011010101",
		340 => "011000000101011010101",
		341 => "011000000101011010101",
		342 => "011010000100001010010",
		343 => "011010000100001010010",
		344 => "011010000100001010010",
		345 => "011000000101011010101",
		346 => "011000000101011010101",
		347 => "011000000101011010101",
		348 => "011001011101001010000",
		349 => "011001011101001010000",
		350 => "011001011101001010000",
		351 => "011000000101011010101",
		352 => "011000000101011010101",
		353 => "011000000101011010101",
		354 => "011010000100001010010",
		355 => "011010000100001010010",
		356 => "011010000100001010010",
		357 => "011000000101011010101",
		358 => "011000000101011010101",
		359 => "011000000101011010101",
		360 => "011001011101001010000",
		361 => "011001011101001010000",
		362 => "011001011101001010000",
		363 => "011000000101011010101",
		364 => "011000000101011010101",
		365 => "011000000101011010101",
		366 => "011010000100001010010",
		367 => "011010000100001010010",
		368 => "011010000100001010010",
		369 => "011000000101011010101",
		370 => "011000000101011010101",
		371 => "011000000101011010101",
		372 => "011001011101001010000",
		373 => "011001011101001010000",
		374 => "011001011101001010000",
		375 => "011000000101011010101",
		376 => "011000000101011010101",
		377 => "011000000101011010101",
		378 => "011010000100001010010",
		379 => "011010000100001010010",
		380 => "011010000100001010010",
		381 => "011000000101011010101",
		382 => "011000000101011010101",
		383 => "011000000101011010101",
		384 => "111011010100001010011",
		385 => "111011010100001010011",
		386 => "111011010100001010011",
		387 => "011000001101100010011",
		388 => "011000001101100010011",
		389 => "011000001101100010011",
		390 => "111011010100001010011",
		391 => "111011010100001010011",
		392 => "111011010100001010011",
		393 => "011000001101100010011",
		394 => "011000001101100010011",
		395 => "011000001101100010011",
		396 => "111011010100001010011",
		397 => "111011010100001010011",
		398 => "111011010100001010011",
		399 => "011000001101100010011",
		400 => "011000001101100010011",
		401 => "011000001101100010011",
		402 => "111011010100001010011",
		403 => "111011010100001010011",
		404 => "111011010100001010011",
		405 => "011000001101100010011",
		406 => "011000001101100010011",
		407 => "011000001101100010011",
		408 => "111011010100001010011",
		409 => "111011010100001010011",
		410 => "111011010100001010011",
		411 => "011000001101100010011",
		412 => "011000001101100010011",
		413 => "011000001101100010011",
		414 => "111011010100001010011",
		415 => "111011010100001010011",
		416 => "111011010100001010011",
		417 => "011000001101100010011",
		418 => "011000001101100010011",
		419 => "011000001101100010011",
		420 => "111011010100001010011",
		421 => "111011010100001010011",
		422 => "111011010100001010011",
		423 => "011000001101100010011",
		424 => "011000001101100010011",
		425 => "011000001101100010011",
		426 => "111011010100001010011",
		427 => "111011010100001010011",
		428 => "111011010100001010011",
		429 => "011000001101100010011",
		430 => "011000001101100010011",
		431 => "011000001101100010011",
		432 => "111011010100001010011",
		433 => "111011010100001010011",
		434 => "111011010100001010011",
		435 => "011000001101100010011",
		436 => "011000001101100010011",
		437 => "011000001101100010011",
		438 => "111011010100001010011",
		439 => "111011010100001010011",
		440 => "111011010100001010011",
		441 => "011000001101100010011",
		442 => "011000001101100010011",
		443 => "011000001101100010011",
		444 => "111011010100001010011",
		445 => "111011010100001010011",
		446 => "111011010100001010011",
		447 => "011000001101100010011",
		448 => "011000001101100010011",
		449 => "011000001101100010011",
		450 => "111011010100001010011",
		451 => "111011010100001010011",
		452 => "111011010100001010011",
		453 => "011000001101100010011",
		454 => "011000001101100010011",
		455 => "011000001101100010011",
		456 => "111011010100001010011",
		457 => "111011010100001010011",
		458 => "111011010100001010011",
		459 => "011000001101100010011",
		460 => "011000001101100010011",
		461 => "011000001101100010011",
		462 => "111011010100001010011",
		463 => "111011010100001010011",
		464 => "111011010100001010011",
		465 => "011000001101100010011",
		466 => "011000001101100010011",
		467 => "011000001101100010011",
		468 => "111011010100001010011",
		469 => "111011010100001010011",
		470 => "111011010100001010011",
		471 => "011000001101100010011",
		472 => "011000001101100010011",
		473 => "011000001101100010011",
		474 => "111011010100001010011",
		475 => "111011010100001010011",
		476 => "111011010100001010011",
		477 => "011000001101100010011",
		478 => "011000001101100010011",
		479 => "011000001101100010011",
		480 => "011011000100001110011",
		481 => "011011000100001110011",
		482 => "011011000100001110011",
		483 => "011011000100001110011",
		484 => "011011000100001110011",
		485 => "011011000100001110011",
		486 => "011011000100001110011",
		487 => "011011000100001110011",
		488 => "011011000100001110011",
		489 => "011011000100001110011",
		490 => "011011000100001110011",
		491 => "011011000100001110011",
		492 => "011011000100001110011",
		493 => "011011000100001110011",
		494 => "011011000100001110011",
		495 => "011011000100001110011",
		496 => "011011000100001110011",
		497 => "011011000100001110011",
		498 => "011011000100001110011",
		499 => "011011000100001110011",
		500 => "011011000100001110011",
		501 => "011011000100001110011",
		502 => "011011000100001110011",
		503 => "011011000100001110011",
		504 => "011011000100001110011",
		505 => "011011000100001110011",
		506 => "011011000100001110011",
		507 => "011011000100001110011",
		508 => "011011000100001110011",
		509 => "011011000100001110011",
		510 => "011011000100001110011",
		511 => "011011000100001110011",
		512 => "011011000100001110011",
		513 => "011011000100001110011",
		514 => "011011000100001110011",
		515 => "011011000100001110011",
		516 => "011011000100001110011",
		517 => "011011000100001110011",
		518 => "011011000100001110011",
		519 => "011011000100001110011",
		520 => "011011000100001110011",
		521 => "011011000100001110011",
		522 => "011011000100001110011",
		523 => "011011000100001110011",
		524 => "011011000100001110011",
		525 => "011011000100001110011",
		526 => "011011000100001110011",
		527 => "011011000100001110011",
		528 => "011011000100001110011",
		529 => "011011000100001110011",
		530 => "011011000100001110011",
		531 => "011011000100001110011",
		532 => "011011000100001110011",
		533 => "011011000100001110011",
		534 => "011011000100001110011",
		535 => "011011000100001110011",
		536 => "011011000100001110011",
		537 => "011011000100001110011",
		538 => "011011000100001110011",
		539 => "011011000100001110011",
		540 => "011011000100001110011",
		541 => "011011000100001110011",
		542 => "011011000100001110011",
		543 => "011011000100001110011",
		544 => "011011000100001110011",
		545 => "011011000100001110011",
		546 => "011011000100001110011",
		547 => "011011000100001110011",
		548 => "011011000100001110011",
		549 => "011011000100001110011",
		550 => "011011000100001110011",
		551 => "011011000100001110011",
		552 => "011011000100001110011",
		553 => "011011000100001110011",
		554 => "011011000100001110011",
		555 => "011011000100001110011",
		556 => "011011000100001110011",
		557 => "011011000100001110011",
		558 => "011011000100001110011",
		559 => "011011000100001110011",
		560 => "011011000100001110011",
		561 => "011011000100001110011",
		562 => "011011000100001110011",
		563 => "011011000100001110011",
		564 => "011011000100001110011",
		565 => "011011000100001110011",
		566 => "011011000100001110011",
		567 => "011011000100001110011",
		568 => "011011000100001110011",
		569 => "011011000100001110011",
		570 => "011011000100001110011",
		571 => "011011000100001110011",
		572 => "011011000100001110011",
		573 => "011011000100001110011",
		574 => "011011000100001110011",
		575 => "011011000100001110011",
		576 => "011000101100100010101",
		577 => "011000101100100010101",
		578 => "011000101100100010101",
		579 => "011000101100100010101",
		580 => "011000101100100010101",
		581 => "011000101100100010101",
		582 => "011000101100100010101",
		583 => "011000101100100010101",
		584 => "011000101100100010101",
		585 => "011000101100100010101",
		586 => "011000101100100010101",
		587 => "011000101100100010101",
		588 => "011000101100100010101",
		589 => "011000101100100010101",
		590 => "011000101100100010101",
		591 => "011000101100100010101",
		592 => "011000101100100010101",
		593 => "011000101100100010101",
		594 => "011000101100100010101",
		595 => "011000101100100010101",
		596 => "011000101100100010101",
		597 => "011000101100100010101",
		598 => "011000101100100010101",
		599 => "011000101100100010101",
		600 => "011000101100100010101",
		601 => "011000101100100010101",
		602 => "011000101100100010101",
		603 => "011000101100100010101",
		604 => "011000101100100010101",
		605 => "011000101100100010101",
		606 => "011000101100100010101",
		607 => "011000101100100010101",
		608 => "011000101100100010101",
		609 => "011000101100100010101",
		610 => "011000101100100010101",
		611 => "011000101100100010101",
		612 => "011000101100100010101",
		613 => "011000101100100010101",
		614 => "011000101100100010101",
		615 => "011000101100100010101",
		616 => "011000101100100010101",
		617 => "011000101100100010101",
		618 => "011000101100100010101",
		619 => "011000101100100010101",
		620 => "011000101100100010101",
		621 => "011000101100100010101",
		622 => "011000101100100010101",
		623 => "011000101100100010101",
		624 => "011000101100100010101",
		625 => "011000101100100010101",
		626 => "011000101100100010101",
		627 => "011000101100100010101",
		628 => "011000101100100010101",
		629 => "011000101100100010101",
		630 => "011000101100100010101",
		631 => "011000101100100010101",
		632 => "011000101100100010101",
		633 => "011000101100100010101",
		634 => "011000101100100010101",
		635 => "011000101100100010101",
		636 => "011000101100100010101",
		637 => "011000101100100010101",
		638 => "011000101100100010101",
		639 => "011000101100100010101",
		640 => "011000101100100010101",
		641 => "011000101100100010101",
		642 => "011000101100100010101",
		643 => "011000101100100010101",
		644 => "011000101100100010101",
		645 => "011000101100100010101",
		646 => "011000101100100010101",
		647 => "011000101100100010101",
		648 => "011000101100100010101",
		649 => "011000101100100010101",
		650 => "011000101100100010101",
		651 => "011000101100100010101",
		652 => "011000101100100010101",
		653 => "011000101100100010101",
		654 => "011000101100100010101",
		655 => "011000101100100010101",
		656 => "011000101100100010101",
		657 => "011000101100100010101",
		658 => "011000101100100010101",
		659 => "011000101100100010101",
		660 => "011000101100100010101",
		661 => "011000101100100010101",
		662 => "011000101100100010101",
		663 => "011000101100100010101",
		664 => "011000101100100010101",
		665 => "011000101100100010101",
		666 => "011000101100100010101",
		667 => "011000101100100010101",
		668 => "011000101100100010101",
		669 => "011000101100100010101",
		670 => "011000101100100010101",
		671 => "011000101100100010101",
		672 => "011000101100100110010",
		673 => "011000101100100110010",
		674 => "011000101100100110010",
		675 => "011000101100100110010",
		676 => "011000101100100110010",
		677 => "011000101100100110010",
		678 => "011000101100100110010",
		679 => "011000101100100110010",
		680 => "011000101100100110010",
		681 => "011000101100100110010",
		682 => "011000101100100110010",
		683 => "011000101100100110010",
		684 => "011000101100100110010",
		685 => "011000101100100110010",
		686 => "011000101100100110010",
		687 => "011000101100100110010",
		688 => "011000101100100110010",
		689 => "011000101100100110010",
		690 => "011000101100100110010",
		691 => "011000101100100110010",
		692 => "011000101100100110010",
		693 => "011000101100100110010",
		694 => "011000101100100110010",
		695 => "011000101100100110010",
		696 => "011000101100100110010",
		697 => "011000101100100110010",
		698 => "011000101100100110010",
		699 => "011000101100100110010",
		700 => "011000101100100110010",
		701 => "011000101100100110010",
		702 => "011000101100100110010",
		703 => "011000101100100110010",
		704 => "011000101100100110010",
		705 => "011000101100100110010",
		706 => "011000101100100110010",
		707 => "011000101100100110010",
		708 => "011000101100100110010",
		709 => "011000101100100110010",
		710 => "011000101100100110010",
		711 => "011000101100100110010",
		712 => "011000101100100110010",
		713 => "011000101100100110010",
		714 => "011000101100100110010",
		715 => "011000101100100110010",
		716 => "011000101100100110010",
		717 => "011000101100100110010",
		718 => "011000101100100110010",
		719 => "011000101100100110010",
		720 => "011000101100100110010",
		721 => "011000101100100110010",
		722 => "011000101100100110010",
		723 => "011000101100100110010",
		724 => "011000101100100110010",
		725 => "011000101100100110010",
		726 => "011000101100100110010",
		727 => "011000101100100110010",
		728 => "011000101100100110010",
		729 => "011000101100100110010",
		730 => "011000101100100110010",
		731 => "011000101100100110010",
		732 => "011000101100100110010",
		733 => "011000101100100110010",
		734 => "011000101100100110010",
		735 => "011000101100100110010",
		736 => "011000101100100110010",
		737 => "011000101100100110010",
		738 => "011000101100100110010",
		739 => "011000101100100110010",
		740 => "011000101100100110010",
		741 => "011000101100100110010",
		742 => "011000101100100110010",
		743 => "011000101100100110010",
		744 => "011000101100100110010",
		745 => "011000101100100110010",
		746 => "011000101100100110010",
		747 => "011000101100100110010",
		748 => "011000101100100110010",
		749 => "011000101100100110010",
		750 => "011000101100100110010",
		751 => "011000101100100110010",
		752 => "011000101100100110010",
		753 => "011000101100100110010",
		754 => "011000101100100110010",
		755 => "011000101100100110010",
		756 => "011000101100100110010",
		757 => "011000101100100110010",
		758 => "011000101100100110010",
		759 => "011000101100100110010",
		760 => "011000101100100110010",
		761 => "011000101100100110010",
		762 => "011000101100100110010",
		763 => "011000101100100110010",
		764 => "011000101100100110010",
		765 => "011000101100100110010",
		766 => "011000101100100110010",
		767 => "011000101100100110010",
		768 => "111000010100001010000",
		769 => "111000010100001010000",
		770 => "111000010100001010000",
		771 => "111000010100001010000",
		772 => "111000010100001010000",
		773 => "111000010100001010000",
		774 => "111000010100001010000",
		775 => "111000010100001010000",
		776 => "111000010100001010000",
		777 => "111000010100001010000",
		778 => "111000010100001010000",
		779 => "111000010100001010000",
		780 => "111000010100001010000",
		781 => "111000010100001010000",
		782 => "111000010100001010000",
		783 => "111000010100001010000",
		784 => "111000010100001010000",
		785 => "111000010100001010000",
		786 => "111000010100001010000",
		787 => "111000010100001010000",
		788 => "111000010100001010000",
		789 => "111000010100001010000",
		790 => "111000010100001010000",
		791 => "111000010100001010000",
		792 => "111000010100001010000",
		793 => "111000010100001010000",
		794 => "111000010100001010000",
		795 => "111000010100001010000",
		796 => "111000010100001010000",
		797 => "111000010100001010000",
		798 => "111000010100001010000",
		799 => "111000010100001010000",
		800 => "111000010100001010000",
		801 => "111000010100001010000",
		802 => "111000010100001010000",
		803 => "111000010100001010000",
		804 => "111000010100001010000",
		805 => "111000010100001010000",
		806 => "111000010100001010000",
		807 => "111000010100001010000",
		808 => "111000010100001010000",
		809 => "111000010100001010000",
		810 => "111000010100001010000",
		811 => "111000010100001010000",
		812 => "111000010100001010000",
		813 => "111000010100001010000",
		814 => "111000010100001010000",
		815 => "111000010100001010000",
		816 => "111000010100001010000",
		817 => "111000010100001010000",
		818 => "111000010100001010000",
		819 => "111000010100001010000",
		820 => "111000010100001010000",
		821 => "111000010100001010000",
		822 => "111000010100001010000",
		823 => "111000010100001010000",
		824 => "111000010100001010000",
		825 => "111000010100001010000",
		826 => "111000010100001010000",
		827 => "111000010100001010000",
		828 => "111000010100001010000",
		829 => "111000010100001010000",
		830 => "111000010100001010000",
		831 => "111000010100001010000",
		832 => "111000010100001010000",
		833 => "111000010100001010000",
		834 => "111000010100001010000",
		835 => "111000010100001010000",
		836 => "111000010100001010000",
		837 => "111000010100001010000",
		838 => "111000010100001010000",
		839 => "111000010100001010000",
		840 => "111000010100001010000",
		841 => "111000010100001010000",
		842 => "111000010100001010000",
		843 => "111000010100001010000",
		844 => "111000010100001010000",
		845 => "111000010100001010000",
		846 => "111000010100001010000",
		847 => "111000010100001010000",
		848 => "111000010100001010000",
		849 => "111000010100001010000",
		850 => "111000010100001010000",
		851 => "111000010100001010000",
		852 => "111000010100001010000",
		853 => "111000010100001010000",
		854 => "111000010100001010000",
		855 => "111000010100001010000",
		856 => "111000010100001010000",
		857 => "111000010100001010000",
		858 => "111000010100001010000",
		859 => "111000010100001010000",
		860 => "111000010100001010000",
		861 => "111000010100001010000",
		862 => "111000010100001010000",
		863 => "111000010100001010000");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;