library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT1024p_6 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT1024p_6;

architecture Behavioral of ROMFFT1024p_6 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 7 
	constant ROM_tb : ROM := (
		0 => "011100001110011010000",
		1 => "011100001110011010000",
		2 => "011100001110011010000",
		3 => "011011100101001110000",
		4 => "011011100101001110000",
		5 => "011011100101001110000",
		6 => "001001111100001010111",
		7 => "001001111100001010111",
		8 => "001001111100001010111",
		9 => "001010011100001010111",
		10 => "001010011100001010111",
		11 => "001010011100001010111",
		12 => "001001011100001010110",
		13 => "001001011100001010110",
		14 => "001001011100001010110",
		15 => "001001111100001010101",
		16 => "001001111100001010101",
		17 => "001001111100001010101",
		18 => "011000111100111010000",
		19 => "011000111100111010000",
		20 => "011000111100111010000",
		21 => "011000110100001010010",
		22 => "011000110100001010010",
		23 => "011000110100001010010",
		24 => "001000011100111010001",
		25 => "001000011100111010001",
		26 => "001000011100111010001",
		27 => "001011011100001010011",
		28 => "001011011100001010011",
		29 => "001011011100001010011",
		30 => "011000111100111010000",
		31 => "011000111100111010000",
		32 => "011000111100111010000",
		33 => "001000100100111110000",
		34 => "001000100100111110000",
		35 => "001000100100111110000",
		36 => "011000000100111010000",
		37 => "011000000100111010000",
		38 => "011000000100111010000",
		39 => "001000111100011110011",
		40 => "001000111100011110011",
		41 => "001000111100011110011",
		42 => "011001100100001110000",
		43 => "011001100100001110000",
		44 => "011001100100001110000",
		45 => "011000011100111010000",
		46 => "011000011100111010000",
		47 => "011000011100111010000",
		48 => "011000000100111010010",
		49 => "011000000100111010010",
		50 => "011000000100111010010",
		51 => "011000001100101010101",
		52 => "011000001100101010101",
		53 => "011000001100101010101",
		54 => "011000000101101010011",
		55 => "011000000101101010011",
		56 => "011000000101101010011",
		57 => "011001111100001010011",
		58 => "011001111100001010011",
		59 => "011001111100001010011",
		60 => "011000000101001010001",
		61 => "011000000101001010001",
		62 => "011000000101001010001",
		63 => "011000000101011010010",
		64 => "011000000101011010010",
		65 => "011000000101011010010",
		66 => "111000011101011010011",
		67 => "111000011101011010011",
		68 => "111000011101011010011",
		69 => "011001100100001110010",
		70 => "011001100100001110010",
		71 => "011001100100001110010",
		72 => "001000011100101110011",
		73 => "001000011100101110011",
		74 => "001000011100101110011",
		75 => "011010100100001110100",
		76 => "011010100100001110100",
		77 => "011010100100001110100",
		78 => "011000000101011010111",
		79 => "011000000101011010111",
		80 => "011000000101011010111",
		81 => "001010111100001010101",
		82 => "001010111100001010101",
		83 => "001010111100001010101",
		84 => "011000000101111010011",
		85 => "011000000101111010011",
		86 => "011000000101111010011",
		87 => "011011011101111010000",
		88 => "011011011101111010000",
		89 => "011011011101111010000",
		90 => "011000001100110110110",
		91 => "011000001100110110110",
		92 => "011000001100110110110",
		93 => "001000011101101011011",
		94 => "001000011101101011011",
		95 => "001000011101101011011",
		96 => "011011101110001010000",
		97 => "011011101110001010000",
		98 => "011011101110001010000",
		99 => "001010011100001010111",
		100 => "001010011100001010111",
		101 => "001010011100001010111",
		102 => "001001100101101110000",
		103 => "001001100101101110000",
		104 => "001001100101101110000",
		105 => "011010100100001010010",
		106 => "011010100100001010010",
		107 => "011010100100001010010",
		108 => "011000001101100010011",
		109 => "011000001101100010011",
		110 => "011000001101100010011",
		111 => "001001011100001010100",
		112 => "001001011100001010100",
		113 => "001001011100001010100",
		114 => "011000001100101010110",
		115 => "011000001100101010110",
		116 => "011000001100101010110",
		117 => "011000011100111010000",
		118 => "011000011100111010000",
		119 => "011000011100111010000",
		120 => "011000101100101010100",
		121 => "011000101100101010100",
		122 => "011000101100101010100",
		123 => "001001111100011110010",
		124 => "001001111100011110010",
		125 => "001001111100011110010",
		126 => "011000000100111010001",
		127 => "011000000100111010001",
		128 => "011000000100111010001",
		129 => "001000110100001010011",
		130 => "001000110100001010011",
		131 => "001000110100001010011",
		132 => "011000000101011010010",
		133 => "011000000101011010010",
		134 => "011000000101011010010",
		135 => "011000000101011010010",
		136 => "011000000101011010010",
		137 => "011000000101011010010",
		138 => "001001111110001010000",
		139 => "001001111110001010000",
		140 => "001001111110001010000",
		141 => "011000000110111010101",
		142 => "011000000110111010101",
		143 => "011000000110111010101",
		144 => "001000011110001010110",
		145 => "001000011110001010110",
		146 => "001000011110001010110",
		147 => "001000011101101010011",
		148 => "001000011101101010011",
		149 => "001000011101101010011",
		150 => "001000010100111010110",
		151 => "001000010100111010110",
		152 => "001000010100111010110",
		153 => "011010100100001010010",
		154 => "011010100100001010010",
		155 => "011010100100001010010",
		156 => "011000001101100010011",
		157 => "011000001101100010011",
		158 => "011000001101100010011",
		159 => "011010000100001010010",
		160 => "011010000100001010010",
		161 => "011010000100001010010",
		162 => "001000111100011110011",
		163 => "001000111100011110011",
		164 => "001000111100011110011",
		165 => "011001000100001110100",
		166 => "011001000100001110100",
		167 => "011001000100001110100",
		168 => "011001000100001110100",
		169 => "011001000100001110100",
		170 => "011001000100001110100",
		171 => "011001000100001010011",
		172 => "011001000100001010011",
		173 => "011001000100001010011",
		174 => "011000000100111010001",
		175 => "011000000100111010001",
		176 => "011000000100111010001",
		177 => "011000101100100110100",
		178 => "011000101100100110100",
		179 => "011000101100100110100",
		180 => "011000000101011010010",
		181 => "011000000101011010010",
		182 => "011000000101011010010",
		183 => "001001011101011010000",
		184 => "001001011101011010000",
		185 => "001001011101011010000",
		186 => "001001111110001010000",
		187 => "001001111110001010000",
		188 => "001001111110001010000",
		189 => "001000011110101010111",
		190 => "001000011110101010111",
		191 => "001000011110101010111",
		192 => "011000000101110011001",
		193 => "011000000101110011001",
		194 => "011000000101110011001",
		195 => "001001111100001010101",
		196 => "001001111100001010101",
		197 => "001001111100001010101",
		198 => "001011011100001010111",
		199 => "001011011100001010111",
		200 => "001011011100001010111",
		201 => "011001011100111010000",
		202 => "011001011100111010000",
		203 => "011001011100111010000",
		204 => "011000000101101010011",
		205 => "011000000101101010011",
		206 => "011000000101101010011",
		207 => "011000001101110010011",
		208 => "011000001101110010011",
		209 => "011000001101110010011",
		210 => "011000001110100010101",
		211 => "011000001110100010101",
		212 => "011000001110100010101",
		213 => "011000000110011010100",
		214 => "011000000110011010100",
		215 => "011000000110011010100",
		216 => "011000000101110011001",
		217 => "011000000101110011001",
		218 => "011000000101110011001",
		219 => "001000011101011010010",
		220 => "001000011101011010010",
		221 => "001000011101011010010",
		222 => "011000111100111010000",
		223 => "011000111100111010000",
		224 => "011000111100111010000",
		225 => "011001100100001010010",
		226 => "011001100100001010010",
		227 => "011001100100001010010",
		228 => "011000000101101010011",
		229 => "011000000101101010011",
		230 => "011000000101101010011",
		231 => "011000001101110010011",
		232 => "011000001101110010011",
		233 => "011000001101110010011",
		234 => "011000001110100010101",
		235 => "011000001110100010101",
		236 => "011000001110100010101",
		237 => "001010011110011010000",
		238 => "001010011110011010000",
		239 => "001010011110011010000",
		240 => "011000000101110011001",
		241 => "011000000101110011001",
		242 => "011000000101110011001",
		243 => "001001111100001010101",
		244 => "001001111100001010101",
		245 => "001001111100001010101",
		246 => "001011011100001010111",
		247 => "001011011100001010111",
		248 => "001011011100001010111",
		249 => "011001011100111010000",
		250 => "011001011100111010000",
		251 => "011001011100111010000",
		252 => "011000000101101010011",
		253 => "011000000101101010011",
		254 => "011000000101101010011",
		255 => "011000001101110010011",
		256 => "011000001101110010011",
		257 => "011000001101110010011",
		258 => "011000001110100010101",
		259 => "011000001110100010101",
		260 => "011000001110100010101",
		261 => "011000000110011010100",
		262 => "011000000110011010100",
		263 => "011000000110011010100",
		264 => "011000000101110011001",
		265 => "011000000101110011001",
		266 => "011000000101110011001",
		267 => "001000011101011010010",
		268 => "001000011101011010010",
		269 => "001000011101011010010",
		270 => "011000111100111010000",
		271 => "011000111100111010000",
		272 => "011000111100111010000",
		273 => "011001100100001010010",
		274 => "011001100100001010010",
		275 => "011001100100001010010",
		276 => "011000000101101010011",
		277 => "011000000101101010011",
		278 => "011000000101101010011",
		279 => "011000001101110010011",
		280 => "011000001101110010011",
		281 => "011000001101110010011",
		282 => "011000001110100010101",
		283 => "011000001110100010101",
		284 => "011000001110100010101",
		285 => "001010011110011010000",
		286 => "001010011110011010000",
		287 => "001010011110011010000",
		288 => "001010111100001010101",
		289 => "001010111100001010101",
		290 => "001010111100001010101",
		291 => "001000111100011110011",
		292 => "001000111100011110011",
		293 => "001000111100011110011",
		294 => "011001011100001010100",
		295 => "011001011100001010100",
		296 => "011001011100001010100",
		297 => "011011100100001110011",
		298 => "011011100100001110011",
		299 => "011011100100001110011",
		300 => "011010100100001010101",
		301 => "011010100100001010101",
		302 => "011010100100001010101",
		303 => "001000100100111010001",
		304 => "001000100100111010001",
		305 => "001000100100111010001",
		306 => "011010000100001110010",
		307 => "011010000100001110010",
		308 => "011010000100001110010",
		309 => "011000000101111010011",
		310 => "011000000101111010011",
		311 => "011000000101111010011",
		312 => "001010111100001010101",
		313 => "001010111100001010101",
		314 => "001010111100001010101",
		315 => "001000111100011110011",
		316 => "001000111100011110011",
		317 => "001000111100011110011",
		318 => "011001011100001010100",
		319 => "011001011100001010100",
		320 => "011001011100001010100",
		321 => "011011100100001110011",
		322 => "011011100100001110011",
		323 => "011011100100001110011",
		324 => "011010100100001010101",
		325 => "011010100100001010101",
		326 => "011010100100001010101",
		327 => "001000100100111010001",
		328 => "001000100100111010001",
		329 => "001000100100111010001",
		330 => "011010000100001110010",
		331 => "011010000100001110010",
		332 => "011010000100001110010",
		333 => "011000000101111010011",
		334 => "011000000101111010011",
		335 => "011000000101111010011",
		336 => "001010111100001010101",
		337 => "001010111100001010101",
		338 => "001010111100001010101",
		339 => "001000111100011110011",
		340 => "001000111100011110011",
		341 => "001000111100011110011",
		342 => "011001011100001010100",
		343 => "011001011100001010100",
		344 => "011001011100001010100",
		345 => "011011100100001110011",
		346 => "011011100100001110011",
		347 => "011011100100001110011",
		348 => "011010100100001010101",
		349 => "011010100100001010101",
		350 => "011010100100001010101",
		351 => "001000100100111010001",
		352 => "001000100100111010001",
		353 => "001000100100111010001",
		354 => "011010000100001110010",
		355 => "011010000100001110010",
		356 => "011010000100001110010",
		357 => "011000000101111010011",
		358 => "011000000101111010011",
		359 => "011000000101111010011",
		360 => "001010111100001010101",
		361 => "001010111100001010101",
		362 => "001010111100001010101",
		363 => "001000111100011110011",
		364 => "001000111100011110011",
		365 => "001000111100011110011",
		366 => "011001011100001010100",
		367 => "011001011100001010100",
		368 => "011001011100001010100",
		369 => "011011100100001110011",
		370 => "011011100100001110011",
		371 => "011011100100001110011",
		372 => "011010100100001010101",
		373 => "011010100100001010101",
		374 => "011010100100001010101",
		375 => "001000100100111010001",
		376 => "001000100100111010001",
		377 => "001000100100111010001",
		378 => "011010000100001110010",
		379 => "011010000100001110010",
		380 => "011010000100001110010",
		381 => "011000000101111010011",
		382 => "011000000101111010011",
		383 => "011000000101111010011",
		384 => "011000001101100010011",
		385 => "011000001101100010011",
		386 => "011000001101100010011",
		387 => "011010100100001010100",
		388 => "011010100100001010100",
		389 => "011010100100001010100",
		390 => "011000001101100010011",
		391 => "011000001101100010011",
		392 => "011000001101100010011",
		393 => "011010100100001010100",
		394 => "011010100100001010100",
		395 => "011010100100001010100",
		396 => "011000001101100010011",
		397 => "011000001101100010011",
		398 => "011000001101100010011",
		399 => "011010100100001010100",
		400 => "011010100100001010100",
		401 => "011010100100001010100",
		402 => "011000001101100010011",
		403 => "011000001101100010011",
		404 => "011000001101100010011",
		405 => "011010100100001010100",
		406 => "011010100100001010100",
		407 => "011010100100001010100",
		408 => "011000001101100010011",
		409 => "011000001101100010011",
		410 => "011000001101100010011",
		411 => "011010100100001010100",
		412 => "011010100100001010100",
		413 => "011010100100001010100",
		414 => "011000001101100010011",
		415 => "011000001101100010011",
		416 => "011000001101100010011",
		417 => "011010100100001010100",
		418 => "011010100100001010100",
		419 => "011010100100001010100",
		420 => "011000001101100010011",
		421 => "011000001101100010011",
		422 => "011000001101100010011",
		423 => "011010100100001010100",
		424 => "011010100100001010100",
		425 => "011010100100001010100",
		426 => "011000001101100010011",
		427 => "011000001101100010011",
		428 => "011000001101100010011",
		429 => "011010100100001010100",
		430 => "011010100100001010100",
		431 => "011010100100001010100",
		432 => "011000001101100010011",
		433 => "011000001101100010011",
		434 => "011000001101100010011",
		435 => "011010100100001010100",
		436 => "011010100100001010100",
		437 => "011010100100001010100",
		438 => "011000001101100010011",
		439 => "011000001101100010011",
		440 => "011000001101100010011",
		441 => "011010100100001010100",
		442 => "011010100100001010100",
		443 => "011010100100001010100",
		444 => "011000001101100010011",
		445 => "011000001101100010011",
		446 => "011000001101100010011",
		447 => "011010100100001010100",
		448 => "011010100100001010100",
		449 => "011010100100001010100",
		450 => "011000001101100010011",
		451 => "011000001101100010011",
		452 => "011000001101100010011",
		453 => "011010100100001010100",
		454 => "011010100100001010100",
		455 => "011010100100001010100",
		456 => "011000001101100010011",
		457 => "011000001101100010011",
		458 => "011000001101100010011",
		459 => "011010100100001010100",
		460 => "011010100100001010100",
		461 => "011010100100001010100",
		462 => "011000001101100010011",
		463 => "011000001101100010011",
		464 => "011000001101100010011",
		465 => "011010100100001010100",
		466 => "011010100100001010100",
		467 => "011010100100001010100",
		468 => "011000001101100010011",
		469 => "011000001101100010011",
		470 => "011000001101100010011",
		471 => "011010100100001010100",
		472 => "011010100100001010100",
		473 => "011010100100001010100",
		474 => "011000001101100010011",
		475 => "011000001101100010011",
		476 => "011000001101100010011",
		477 => "011010100100001010100",
		478 => "011010100100001010100",
		479 => "011010100100001010100",
		480 => "011001100100001110001",
		481 => "011001100100001110001",
		482 => "011001100100001110001",
		483 => "001000111100111010000",
		484 => "001000111100111010000",
		485 => "001000111100111010000",
		486 => "011001100100001110001",
		487 => "011001100100001110001",
		488 => "011001100100001110001",
		489 => "001000111100111010000",
		490 => "001000111100111010000",
		491 => "001000111100111010000",
		492 => "011001100100001110001",
		493 => "011001100100001110001",
		494 => "011001100100001110001",
		495 => "001000111100111010000",
		496 => "001000111100111010000",
		497 => "001000111100111010000",
		498 => "011001100100001110001",
		499 => "011001100100001110001",
		500 => "011001100100001110001",
		501 => "001000111100111010000",
		502 => "001000111100111010000",
		503 => "001000111100111010000",
		504 => "011001100100001110001",
		505 => "011001100100001110001",
		506 => "011001100100001110001",
		507 => "001000111100111010000",
		508 => "001000111100111010000",
		509 => "001000111100111010000",
		510 => "011001100100001110001",
		511 => "011001100100001110001",
		512 => "011001100100001110001",
		513 => "001000111100111010000",
		514 => "001000111100111010000",
		515 => "001000111100111010000",
		516 => "011001100100001110001",
		517 => "011001100100001110001",
		518 => "011001100100001110001",
		519 => "001000111100111010000",
		520 => "001000111100111010000",
		521 => "001000111100111010000",
		522 => "011001100100001110001",
		523 => "011001100100001110001",
		524 => "011001100100001110001",
		525 => "001000111100111010000",
		526 => "001000111100111010000",
		527 => "001000111100111010000",
		528 => "011001100100001110001",
		529 => "011001100100001110001",
		530 => "011001100100001110001",
		531 => "001000111100111010000",
		532 => "001000111100111010000",
		533 => "001000111100111010000",
		534 => "011001100100001110001",
		535 => "011001100100001110001",
		536 => "011001100100001110001",
		537 => "001000111100111010000",
		538 => "001000111100111010000",
		539 => "001000111100111010000",
		540 => "011001100100001110001",
		541 => "011001100100001110001",
		542 => "011001100100001110001",
		543 => "001000111100111010000",
		544 => "001000111100111010000",
		545 => "001000111100111010000",
		546 => "011001100100001110001",
		547 => "011001100100001110001",
		548 => "011001100100001110001",
		549 => "001000111100111010000",
		550 => "001000111100111010000",
		551 => "001000111100111010000",
		552 => "011001100100001110001",
		553 => "011001100100001110001",
		554 => "011001100100001110001",
		555 => "001000111100111010000",
		556 => "001000111100111010000",
		557 => "001000111100111010000",
		558 => "011001100100001110001",
		559 => "011001100100001110001",
		560 => "011001100100001110001",
		561 => "001000111100111010000",
		562 => "001000111100111010000",
		563 => "001000111100111010000",
		564 => "011001100100001110001",
		565 => "011001100100001110001",
		566 => "011001100100001110001",
		567 => "001000111100111010000",
		568 => "001000111100111010000",
		569 => "001000111100111010000",
		570 => "011001100100001110001",
		571 => "011001100100001110001",
		572 => "011001100100001110001",
		573 => "001000111100111010000",
		574 => "001000111100111010000",
		575 => "001000111100111010000",
		576 => "011000101100100010101",
		577 => "011000101100100010101",
		578 => "011000101100100010101",
		579 => "011000101100100010101",
		580 => "011000101100100010101",
		581 => "011000101100100010101",
		582 => "011000101100100010101",
		583 => "011000101100100010101",
		584 => "011000101100100010101",
		585 => "011000101100100010101",
		586 => "011000101100100010101",
		587 => "011000101100100010101",
		588 => "011000101100100010101",
		589 => "011000101100100010101",
		590 => "011000101100100010101",
		591 => "011000101100100010101",
		592 => "011000101100100010101",
		593 => "011000101100100010101",
		594 => "011000101100100010101",
		595 => "011000101100100010101",
		596 => "011000101100100010101",
		597 => "011000101100100010101",
		598 => "011000101100100010101",
		599 => "011000101100100010101",
		600 => "011000101100100010101",
		601 => "011000101100100010101",
		602 => "011000101100100010101",
		603 => "011000101100100010101",
		604 => "011000101100100010101",
		605 => "011000101100100010101",
		606 => "011000101100100010101",
		607 => "011000101100100010101",
		608 => "011000101100100010101",
		609 => "011000101100100010101",
		610 => "011000101100100010101",
		611 => "011000101100100010101",
		612 => "011000101100100010101",
		613 => "011000101100100010101",
		614 => "011000101100100010101",
		615 => "011000101100100010101",
		616 => "011000101100100010101",
		617 => "011000101100100010101",
		618 => "011000101100100010101",
		619 => "011000101100100010101",
		620 => "011000101100100010101",
		621 => "011000101100100010101",
		622 => "011000101100100010101",
		623 => "011000101100100010101",
		624 => "011000101100100010101",
		625 => "011000101100100010101",
		626 => "011000101100100010101",
		627 => "011000101100100010101",
		628 => "011000101100100010101",
		629 => "011000101100100010101",
		630 => "011000101100100010101",
		631 => "011000101100100010101",
		632 => "011000101100100010101",
		633 => "011000101100100010101",
		634 => "011000101100100010101",
		635 => "011000101100100010101",
		636 => "011000101100100010101",
		637 => "011000101100100010101",
		638 => "011000101100100010101",
		639 => "011000101100100010101",
		640 => "011000101100100010101",
		641 => "011000101100100010101",
		642 => "011000101100100010101",
		643 => "011000101100100010101",
		644 => "011000101100100010101",
		645 => "011000101100100010101",
		646 => "011000101100100010101",
		647 => "011000101100100010101",
		648 => "011000101100100010101",
		649 => "011000101100100010101",
		650 => "011000101100100010101",
		651 => "011000101100100010101",
		652 => "011000101100100010101",
		653 => "011000101100100010101",
		654 => "011000101100100010101",
		655 => "011000101100100010101",
		656 => "011000101100100010101",
		657 => "011000101100100010101",
		658 => "011000101100100010101",
		659 => "011000101100100010101",
		660 => "011000101100100010101",
		661 => "011000101100100010101",
		662 => "011000101100100010101",
		663 => "011000101100100010101",
		664 => "011000101100100010101",
		665 => "011000101100100010101",
		666 => "011000101100100010101",
		667 => "011000101100100010101",
		668 => "011000101100100010101",
		669 => "011000101100100010101",
		670 => "011000101100100010101",
		671 => "011000101100100010101",
		672 => "011000101100100110010",
		673 => "011000101100100110010",
		674 => "011000101100100110010",
		675 => "011000101100100110010",
		676 => "011000101100100110010",
		677 => "011000101100100110010",
		678 => "011000101100100110010",
		679 => "011000101100100110010",
		680 => "011000101100100110010",
		681 => "011000101100100110010",
		682 => "011000101100100110010",
		683 => "011000101100100110010",
		684 => "011000101100100110010",
		685 => "011000101100100110010",
		686 => "011000101100100110010",
		687 => "011000101100100110010",
		688 => "011000101100100110010",
		689 => "011000101100100110010",
		690 => "011000101100100110010",
		691 => "011000101100100110010",
		692 => "011000101100100110010",
		693 => "011000101100100110010",
		694 => "011000101100100110010",
		695 => "011000101100100110010",
		696 => "011000101100100110010",
		697 => "011000101100100110010",
		698 => "011000101100100110010",
		699 => "011000101100100110010",
		700 => "011000101100100110010",
		701 => "011000101100100110010",
		702 => "011000101100100110010",
		703 => "011000101100100110010",
		704 => "011000101100100110010",
		705 => "011000101100100110010",
		706 => "011000101100100110010",
		707 => "011000101100100110010",
		708 => "011000101100100110010",
		709 => "011000101100100110010",
		710 => "011000101100100110010",
		711 => "011000101100100110010",
		712 => "011000101100100110010",
		713 => "011000101100100110010",
		714 => "011000101100100110010",
		715 => "011000101100100110010",
		716 => "011000101100100110010",
		717 => "011000101100100110010",
		718 => "011000101100100110010",
		719 => "011000101100100110010",
		720 => "011000101100100110010",
		721 => "011000101100100110010",
		722 => "011000101100100110010",
		723 => "011000101100100110010",
		724 => "011000101100100110010",
		725 => "011000101100100110010",
		726 => "011000101100100110010",
		727 => "011000101100100110010",
		728 => "011000101100100110010",
		729 => "011000101100100110010",
		730 => "011000101100100110010",
		731 => "011000101100100110010",
		732 => "011000101100100110010",
		733 => "011000101100100110010",
		734 => "011000101100100110010",
		735 => "011000101100100110010",
		736 => "011000101100100110010",
		737 => "011000101100100110010",
		738 => "011000101100100110010",
		739 => "011000101100100110010",
		740 => "011000101100100110010",
		741 => "011000101100100110010",
		742 => "011000101100100110010",
		743 => "011000101100100110010",
		744 => "011000101100100110010",
		745 => "011000101100100110010",
		746 => "011000101100100110010",
		747 => "011000101100100110010",
		748 => "011000101100100110010",
		749 => "011000101100100110010",
		750 => "011000101100100110010",
		751 => "011000101100100110010",
		752 => "011000101100100110010",
		753 => "011000101100100110010",
		754 => "011000101100100110010",
		755 => "011000101100100110010",
		756 => "011000101100100110010",
		757 => "011000101100100110010",
		758 => "011000101100100110010",
		759 => "011000101100100110010",
		760 => "011000101100100110010",
		761 => "011000101100100110010",
		762 => "011000101100100110010",
		763 => "011000101100100110010",
		764 => "011000101100100110010",
		765 => "011000101100100110010",
		766 => "011000101100100110010",
		767 => "011000101100100110010",
		768 => "111000010100001010000",
		769 => "111000010100001010000",
		770 => "111000010100001010000",
		771 => "111000010100001010000",
		772 => "111000010100001010000",
		773 => "111000010100001010000",
		774 => "111000010100001010000",
		775 => "111000010100001010000",
		776 => "111000010100001010000",
		777 => "111000010100001010000",
		778 => "111000010100001010000",
		779 => "111000010100001010000",
		780 => "111000010100001010000",
		781 => "111000010100001010000",
		782 => "111000010100001010000",
		783 => "111000010100001010000",
		784 => "111000010100001010000",
		785 => "111000010100001010000",
		786 => "111000010100001010000",
		787 => "111000010100001010000",
		788 => "111000010100001010000",
		789 => "111000010100001010000",
		790 => "111000010100001010000",
		791 => "111000010100001010000",
		792 => "111000010100001010000",
		793 => "111000010100001010000",
		794 => "111000010100001010000",
		795 => "111000010100001010000",
		796 => "111000010100001010000",
		797 => "111000010100001010000",
		798 => "111000010100001010000",
		799 => "111000010100001010000",
		800 => "111000010100001010000",
		801 => "111000010100001010000",
		802 => "111000010100001010000",
		803 => "111000010100001010000",
		804 => "111000010100001010000",
		805 => "111000010100001010000",
		806 => "111000010100001010000",
		807 => "111000010100001010000",
		808 => "111000010100001010000",
		809 => "111000010100001010000",
		810 => "111000010100001010000",
		811 => "111000010100001010000",
		812 => "111000010100001010000",
		813 => "111000010100001010000",
		814 => "111000010100001010000",
		815 => "111000010100001010000",
		816 => "111000010100001010000",
		817 => "111000010100001010000",
		818 => "111000010100001010000",
		819 => "111000010100001010000",
		820 => "111000010100001010000",
		821 => "111000010100001010000",
		822 => "111000010100001010000",
		823 => "111000010100001010000",
		824 => "111000010100001010000",
		825 => "111000010100001010000",
		826 => "111000010100001010000",
		827 => "111000010100001010000",
		828 => "111000010100001010000",
		829 => "111000010100001010000",
		830 => "111000010100001010000",
		831 => "111000010100001010000",
		832 => "111000010100001010000",
		833 => "111000010100001010000",
		834 => "111000010100001010000",
		835 => "111000010100001010000",
		836 => "111000010100001010000",
		837 => "111000010100001010000",
		838 => "111000010100001010000",
		839 => "111000010100001010000",
		840 => "111000010100001010000",
		841 => "111000010100001010000",
		842 => "111000010100001010000",
		843 => "111000010100001010000",
		844 => "111000010100001010000",
		845 => "111000010100001010000",
		846 => "111000010100001010000",
		847 => "111000010100001010000",
		848 => "111000010100001010000",
		849 => "111000010100001010000",
		850 => "111000010100001010000",
		851 => "111000010100001010000",
		852 => "111000010100001010000",
		853 => "111000010100001010000",
		854 => "111000010100001010000",
		855 => "111000010100001010000",
		856 => "111000010100001010000",
		857 => "111000010100001010000",
		858 => "111000010100001010000",
		859 => "111000010100001010000",
		860 => "111000010100001010000",
		861 => "111000010100001010000",
		862 => "111000010100001010000",
		863 => "111000010100001010000");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;