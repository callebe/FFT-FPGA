library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT8 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT8;

architecture Behavioral of ROMFFT8 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 9 
	constant ROM_tb : ROM := (
		0 => "011000000110011110100",
		1 => "011000000110011110100",
		2 => "011000000110011110100",
		3 => "011000000101110011001",
		4 => "011000000101110011001",
		5 => "011000000101110011001",
		6 => "011000001110100010101",
		7 => "011000001110100010101",
		8 => "011000001110100010101",
		9 => "001001111100001010101",
		10 => "001001111100001010101",
		11 => "001001111100001010101",
		12 => "011000000100111010110",
		13 => "011000000100111010110",
		14 => "011000000100111010110",
		15 => "001011011100001010111",
		16 => "001011011100001010111",
		17 => "001011011100001010111",
		18 => "001001111100001010110",
		19 => "001001111100001010110",
		20 => "001001111100001010110",
		21 => "011001011100111010000",
		22 => "011001011100111010000",
		23 => "011001011100111010000",
		24 => "011001011100001010011",
		25 => "011001011100001010011",
		26 => "011001011100001010011",
		27 => "011000000101101010011",
		28 => "011000000101101010011",
		29 => "011000000101101010011",
		30 => "011000111100001010011",
		31 => "011000111100001010011",
		32 => "011000111100001010011",
		33 => "011000001101110010011",
		34 => "011000001101110010011",
		35 => "011000001101110010011",
		36 => "011000000101011010011",
		37 => "011000000101011010011",
		38 => "011000000101011010011",
		39 => "011000001110100010101",
		40 => "011000001110100010101",
		41 => "011000001110100010101",
		42 => "011000010100111010110",
		43 => "011000010100111010110",
		44 => "011000010100111010110",
		45 => "011000000110011010100",
		46 => "011000000110011010100",
		47 => "011000000110011010100",
		48 => "001010011100001011001",
		49 => "001010011100001011001",
		50 => "001010011100001011001",
		51 => "011000000101110011001",
		52 => "011000000101110011001",
		53 => "011000000101110011001",
		54 => "011000001110100010101",
		55 => "011000001110100010101",
		56 => "011000001110100010101",
		57 => "001000011101011010010",
		58 => "001000011101011010010",
		59 => "001000011101011010010",
		60 => "011000001101110010011",
		61 => "011000001101110010011",
		62 => "011000001101110010011",
		63 => "011000111100111010000",
		64 => "011000111100111010000",
		65 => "011000111100111010000",
		66 => "011011000100001010011",
		67 => "011011000100001010011",
		68 => "011011000100001010011",
		69 => "011001100100001010010",
		70 => "011001100100001010010",
		71 => "011001100100001010010",
		72 => "011001100100001110010",
		73 => "011001100100001110010",
		74 => "011001100100001110010",
		75 => "011000000101101010011",
		76 => "011000000101101010011",
		77 => "011000000101101010011",
		78 => "011001100100001110001",
		79 => "011001100100001110001",
		80 => "011001100100001110001",
		81 => "011000001101110010011",
		82 => "011000001101110010011",
		83 => "011000001101110010011",
		84 => "011010100100001110011",
		85 => "011010100100001110011",
		86 => "011010100100001110011",
		87 => "011000001110100010101",
		88 => "011000001110100010101",
		89 => "011000001110100010101",
		90 => "011000000101110011001",
		91 => "011000000101110011001",
		92 => "011000000101110011001",
		93 => "001010011110011010000",
		94 => "001010011110011010000",
		95 => "001010011110011010000",
		96 => "011000000101111110011",
		97 => "011000000101111110011",
		98 => "011000000101111110011",
		99 => "001010111100001010101",
		100 => "001010111100001010101",
		101 => "001010111100001010101",
		102 => "011001011101001010000",
		103 => "011001011101001010000",
		104 => "011001011101001010000",
		105 => "001000111100011110011",
		106 => "001000111100011110011",
		107 => "001000111100011110011",
		108 => "011000101100111010001",
		109 => "011000101100111010001",
		110 => "011000101100111010001",
		111 => "011001011100001010100",
		112 => "011001011100001010100",
		113 => "011001011100001010100",
		114 => "011000000101011010101",
		115 => "011000000101011010101",
		116 => "011000000101011010101",
		117 => "011011100100001110011",
		118 => "011011100100001110011",
		119 => "011011100100001110011",
		120 => "001001111100001010111",
		121 => "001001111100001010111",
		122 => "001001111100001010111",
		123 => "011010100100001010101",
		124 => "011010100100001010101",
		125 => "011010100100001010101",
		126 => "011010000100001010010",
		127 => "011010000100001010010",
		128 => "011010000100001010010",
		129 => "001000100100111010001",
		130 => "001000100100111010001",
		131 => "001000100100111010001",
		132 => "001000000100101110110",
		133 => "001000000100101110110",
		134 => "001000000100101110110",
		135 => "011010000100001110010",
		136 => "011010000100001110010",
		137 => "011010000100001110010",
		138 => "011000000101011010101",
		139 => "011000000101011010101",
		140 => "011000000101011010101",
		141 => "011000000101111010011",
		142 => "011000000101111010011",
		143 => "011000000101111010011",
		144 => "011000000101111110011",
		145 => "011000000101111110011",
		146 => "011000000101111110011",
		147 => "001010111100001010101",
		148 => "001010111100001010101",
		149 => "001010111100001010101",
		150 => "011001011101001010000",
		151 => "011001011101001010000",
		152 => "011001011101001010000",
		153 => "001000111100011110011",
		154 => "001000111100011110011",
		155 => "001000111100011110011",
		156 => "011000101100111010001",
		157 => "011000101100111010001",
		158 => "011000101100111010001",
		159 => "011001011100001010100",
		160 => "011001011100001010100",
		161 => "011001011100001010100",
		162 => "011000000101011010101",
		163 => "011000000101011010101",
		164 => "011000000101011010101",
		165 => "011011100100001110011",
		166 => "011011100100001110011",
		167 => "011011100100001110011",
		168 => "001001111100001010111",
		169 => "001001111100001010111",
		170 => "001001111100001010111",
		171 => "011010100100001010101",
		172 => "011010100100001010101",
		173 => "011010100100001010101",
		174 => "011010000100001010010",
		175 => "011010000100001010010",
		176 => "011010000100001010010",
		177 => "001000100100111010001",
		178 => "001000100100111010001",
		179 => "001000100100111010001",
		180 => "001000000100101110110",
		181 => "001000000100101110110",
		182 => "001000000100101110110",
		183 => "011010000100001110010",
		184 => "011010000100001110010",
		185 => "011010000100001110010",
		186 => "011000000101011010101",
		187 => "011000000101011010101",
		188 => "011000000101011010101",
		189 => "011000000101111010011",
		190 => "011000000101111010011",
		191 => "011000000101111010011",
		192 => "011010100100001110100",
		193 => "011010100100001110100",
		194 => "011010100100001110100",
		195 => "011000001101100010011",
		196 => "011000001101100010011",
		197 => "011000001101100010011",
		198 => "111011010100001010011",
		199 => "111011010100001010011",
		200 => "111011010100001010011",
		201 => "011010100100001010100",
		202 => "011010100100001010100",
		203 => "011010100100001010100",
		204 => "011010100100001110100",
		205 => "011010100100001110100",
		206 => "011010100100001110100",
		207 => "011000001101100010011",
		208 => "011000001101100010011",
		209 => "011000001101100010011",
		210 => "011000001101100010011",
		211 => "011000001101100010011",
		212 => "011000001101100010011",
		213 => "011010100100001010100",
		214 => "011010100100001010100",
		215 => "011010100100001010100",
		216 => "011010100100001110100",
		217 => "011010100100001110100",
		218 => "011010100100001110100",
		219 => "011000001101100010011",
		220 => "011000001101100010011",
		221 => "011000001101100010011",
		222 => "111011010100001010011",
		223 => "111011010100001010011",
		224 => "111011010100001010011",
		225 => "011010100100001010100",
		226 => "011010100100001010100",
		227 => "011010100100001010100",
		228 => "011010100100001110100",
		229 => "011010100100001110100",
		230 => "011010100100001110100",
		231 => "011000001101100010011",
		232 => "011000001101100010011",
		233 => "011000001101100010011",
		234 => "011000001101100010011",
		235 => "011000001101100010011",
		236 => "011000001101100010011",
		237 => "011010100100001010100",
		238 => "011010100100001010100",
		239 => "011010100100001010100",
		240 => "011010100100001110100",
		241 => "011010100100001110100",
		242 => "011010100100001110100",
		243 => "011000001101100010011",
		244 => "011000001101100010011",
		245 => "011000001101100010011",
		246 => "111011010100001010011",
		247 => "111011010100001010011",
		248 => "111011010100001010011",
		249 => "011010100100001010100",
		250 => "011010100100001010100",
		251 => "011010100100001010100",
		252 => "011010100100001110100",
		253 => "011010100100001110100",
		254 => "011010100100001110100",
		255 => "011000001101100010011",
		256 => "011000001101100010011",
		257 => "011000001101100010011",
		258 => "011000001101100010011",
		259 => "011000001101100010011",
		260 => "011000001101100010011",
		261 => "011010100100001010100",
		262 => "011010100100001010100",
		263 => "011010100100001010100",
		264 => "011010100100001110100",
		265 => "011010100100001110100",
		266 => "011010100100001110100",
		267 => "011000001101100010011",
		268 => "011000001101100010011",
		269 => "011000001101100010011",
		270 => "111011010100001010011",
		271 => "111011010100001010011",
		272 => "111011010100001010011",
		273 => "011010100100001010100",
		274 => "011010100100001010100",
		275 => "011010100100001010100",
		276 => "011010100100001110100",
		277 => "011010100100001110100",
		278 => "011010100100001110100",
		279 => "011000001101100010011",
		280 => "011000001101100010011",
		281 => "011000001101100010011",
		282 => "011000001101100010011",
		283 => "011000001101100010011",
		284 => "011000001101100010011",
		285 => "011010100100001010100",
		286 => "011010100100001010100",
		287 => "011010100100001010100",
		288 => "011001111100001010110",
		289 => "011001111100001010110",
		290 => "011001111100001010110",
		291 => "011001100100001110001",
		292 => "011001100100001110001",
		293 => "011001100100001110001",
		294 => "011011000100001110011",
		295 => "011011000100001110011",
		296 => "011011000100001110011",
		297 => "001000111100111010000",
		298 => "001000111100111010000",
		299 => "001000111100111010000",
		300 => "011001111100001010110",
		301 => "011001111100001010110",
		302 => "011001111100001010110",
		303 => "011001100100001110001",
		304 => "011001100100001110001",
		305 => "011001100100001110001",
		306 => "011011000100001110011",
		307 => "011011000100001110011",
		308 => "011011000100001110011",
		309 => "001000111100111010000",
		310 => "001000111100111010000",
		311 => "001000111100111010000",
		312 => "011001111100001010110",
		313 => "011001111100001010110",
		314 => "011001111100001010110",
		315 => "011001100100001110001",
		316 => "011001100100001110001",
		317 => "011001100100001110001",
		318 => "011011000100001110011",
		319 => "011011000100001110011",
		320 => "011011000100001110011",
		321 => "001000111100111010000",
		322 => "001000111100111010000",
		323 => "001000111100111010000",
		324 => "011001111100001010110",
		325 => "011001111100001010110",
		326 => "011001111100001010110",
		327 => "011001100100001110001",
		328 => "011001100100001110001",
		329 => "011001100100001110001",
		330 => "011011000100001110011",
		331 => "011011000100001110011",
		332 => "011011000100001110011",
		333 => "001000111100111010000",
		334 => "001000111100111010000",
		335 => "001000111100111010000",
		336 => "011001111100001010110",
		337 => "011001111100001010110",
		338 => "011001111100001010110",
		339 => "011001100100001110001",
		340 => "011001100100001110001",
		341 => "011001100100001110001",
		342 => "011011000100001110011",
		343 => "011011000100001110011",
		344 => "011011000100001110011",
		345 => "001000111100111010000",
		346 => "001000111100111010000",
		347 => "001000111100111010000",
		348 => "011001111100001010110",
		349 => "011001111100001010110",
		350 => "011001111100001010110",
		351 => "011001100100001110001",
		352 => "011001100100001110001",
		353 => "011001100100001110001",
		354 => "011011000100001110011",
		355 => "011011000100001110011",
		356 => "011011000100001110011",
		357 => "001000111100111010000",
		358 => "001000111100111010000",
		359 => "001000111100111010000",
		360 => "011001111100001010110",
		361 => "011001111100001010110",
		362 => "011001111100001010110",
		363 => "011001100100001110001",
		364 => "011001100100001110001",
		365 => "011001100100001110001",
		366 => "011011000100001110011",
		367 => "011011000100001110011",
		368 => "011011000100001110011",
		369 => "001000111100111010000",
		370 => "001000111100111010000",
		371 => "001000111100111010000",
		372 => "011001111100001010110",
		373 => "011001111100001010110",
		374 => "011001111100001010110",
		375 => "011001100100001110001",
		376 => "011001100100001110001",
		377 => "011001100100001110001",
		378 => "011011000100001110011",
		379 => "011011000100001110011",
		380 => "011011000100001110011",
		381 => "001000111100111010000",
		382 => "001000111100111010000",
		383 => "001000111100111010000",
		384 => "011000101100100010101",
		385 => "011000101100100010101",
		386 => "011000101100100010101",
		387 => "011000101100100010101",
		388 => "011000101100100010101",
		389 => "011000101100100010101",
		390 => "011000101100100010101",
		391 => "011000101100100010101",
		392 => "011000101100100010101",
		393 => "011000101100100010101",
		394 => "011000101100100010101",
		395 => "011000101100100010101",
		396 => "011000101100100010101",
		397 => "011000101100100010101",
		398 => "011000101100100010101",
		399 => "011000101100100010101",
		400 => "011000101100100010101",
		401 => "011000101100100010101",
		402 => "011000101100100010101",
		403 => "011000101100100010101",
		404 => "011000101100100010101",
		405 => "011000101100100010101",
		406 => "011000101100100010101",
		407 => "011000101100100010101",
		408 => "011000101100100010101",
		409 => "011000101100100010101",
		410 => "011000101100100010101",
		411 => "011000101100100010101",
		412 => "011000101100100010101",
		413 => "011000101100100010101",
		414 => "011000101100100010101",
		415 => "011000101100100010101",
		416 => "011000101100100010101",
		417 => "011000101100100010101",
		418 => "011000101100100010101",
		419 => "011000101100100010101",
		420 => "011000101100100010101",
		421 => "011000101100100010101",
		422 => "011000101100100010101",
		423 => "011000101100100010101",
		424 => "011000101100100010101",
		425 => "011000101100100010101",
		426 => "011000101100100010101",
		427 => "011000101100100010101",
		428 => "011000101100100010101",
		429 => "011000101100100010101",
		430 => "011000101100100010101",
		431 => "011000101100100010101",
		432 => "011000101100100010101",
		433 => "011000101100100010101",
		434 => "011000101100100010101",
		435 => "011000101100100010101",
		436 => "011000101100100010101",
		437 => "011000101100100010101",
		438 => "011000101100100010101",
		439 => "011000101100100010101",
		440 => "011000101100100010101",
		441 => "011000101100100010101",
		442 => "011000101100100010101",
		443 => "011000101100100010101",
		444 => "011000101100100010101",
		445 => "011000101100100010101",
		446 => "011000101100100010101",
		447 => "011000101100100010101",
		448 => "011000101100100010101",
		449 => "011000101100100010101",
		450 => "011000101100100010101",
		451 => "011000101100100010101",
		452 => "011000101100100010101",
		453 => "011000101100100010101",
		454 => "011000101100100010101",
		455 => "011000101100100010101",
		456 => "011000101100100010101",
		457 => "011000101100100010101",
		458 => "011000101100100010101",
		459 => "011000101100100010101",
		460 => "011000101100100010101",
		461 => "011000101100100010101",
		462 => "011000101100100010101",
		463 => "011000101100100010101",
		464 => "011000101100100010101",
		465 => "011000101100100010101",
		466 => "011000101100100010101",
		467 => "011000101100100010101",
		468 => "011000101100100010101",
		469 => "011000101100100010101",
		470 => "011000101100100010101",
		471 => "011000101100100010101",
		472 => "011000101100100010101",
		473 => "011000101100100010101",
		474 => "011000101100100010101",
		475 => "011000101100100010101",
		476 => "011000101100100010101",
		477 => "011000101100100010101",
		478 => "011000101100100010101",
		479 => "011000101100100010101",
		480 => "011000101100100110010",
		481 => "011000101100100110010",
		482 => "011000101100100110010",
		483 => "011000101100100110010",
		484 => "011000101100100110010",
		485 => "011000101100100110010",
		486 => "011000101100100110010",
		487 => "011000101100100110010",
		488 => "011000101100100110010",
		489 => "011000101100100110010",
		490 => "011000101100100110010",
		491 => "011000101100100110010",
		492 => "011000101100100110010",
		493 => "011000101100100110010",
		494 => "011000101100100110010",
		495 => "011000101100100110010",
		496 => "011000101100100110010",
		497 => "011000101100100110010",
		498 => "011000101100100110010",
		499 => "011000101100100110010",
		500 => "011000101100100110010",
		501 => "011000101100100110010",
		502 => "011000101100100110010",
		503 => "011000101100100110010",
		504 => "011000101100100110010",
		505 => "011000101100100110010",
		506 => "011000101100100110010",
		507 => "011000101100100110010",
		508 => "011000101100100110010",
		509 => "011000101100100110010",
		510 => "011000101100100110010",
		511 => "011000101100100110010",
		512 => "011000101100100110010",
		513 => "011000101100100110010",
		514 => "011000101100100110010",
		515 => "011000101100100110010",
		516 => "011000101100100110010",
		517 => "011000101100100110010",
		518 => "011000101100100110010",
		519 => "011000101100100110010",
		520 => "011000101100100110010",
		521 => "011000101100100110010",
		522 => "011000101100100110010",
		523 => "011000101100100110010",
		524 => "011000101100100110010",
		525 => "011000101100100110010",
		526 => "011000101100100110010",
		527 => "011000101100100110010",
		528 => "011000101100100110010",
		529 => "011000101100100110010",
		530 => "011000101100100110010",
		531 => "011000101100100110010",
		532 => "011000101100100110010",
		533 => "011000101100100110010",
		534 => "011000101100100110010",
		535 => "011000101100100110010",
		536 => "011000101100100110010",
		537 => "011000101100100110010",
		538 => "011000101100100110010",
		539 => "011000101100100110010",
		540 => "011000101100100110010",
		541 => "011000101100100110010",
		542 => "011000101100100110010",
		543 => "011000101100100110010",
		544 => "011000101100100110010",
		545 => "011000101100100110010",
		546 => "011000101100100110010",
		547 => "011000101100100110010",
		548 => "011000101100100110010",
		549 => "011000101100100110010",
		550 => "011000101100100110010",
		551 => "011000101100100110010",
		552 => "011000101100100110010",
		553 => "011000101100100110010",
		554 => "011000101100100110010",
		555 => "011000101100100110010",
		556 => "011000101100100110010",
		557 => "011000101100100110010",
		558 => "011000101100100110010",
		559 => "011000101100100110010",
		560 => "011000101100100110010",
		561 => "011000101100100110010",
		562 => "011000101100100110010",
		563 => "011000101100100110010",
		564 => "011000101100100110010",
		565 => "011000101100100110010",
		566 => "011000101100100110010",
		567 => "011000101100100110010",
		568 => "011000101100100110010",
		569 => "011000101100100110010",
		570 => "011000101100100110010",
		571 => "011000101100100110010",
		572 => "011000101100100110010",
		573 => "011000101100100110010",
		574 => "011000101100100110010",
		575 => "011000101100100110010",
		576 => "111000010100001010000",
		577 => "111000010100001010000",
		578 => "111000010100001010000",
		579 => "111000010100001010000",
		580 => "111000010100001010000",
		581 => "111000010100001010000",
		582 => "111000010100001010000",
		583 => "111000010100001010000",
		584 => "111000010100001010000",
		585 => "111000010100001010000",
		586 => "111000010100001010000",
		587 => "111000010100001010000",
		588 => "111000010100001010000",
		589 => "111000010100001010000",
		590 => "111000010100001010000",
		591 => "111000010100001010000",
		592 => "111000010100001010000",
		593 => "111000010100001010000",
		594 => "111000010100001010000",
		595 => "111000010100001010000",
		596 => "111000010100001010000",
		597 => "111000010100001010000",
		598 => "111000010100001010000",
		599 => "111000010100001010000",
		600 => "111000010100001010000",
		601 => "111000010100001010000",
		602 => "111000010100001010000",
		603 => "111000010100001010000",
		604 => "111000010100001010000",
		605 => "111000010100001010000",
		606 => "111000010100001010000",
		607 => "111000010100001010000",
		608 => "111000010100001010000",
		609 => "111000010100001010000",
		610 => "111000010100001010000",
		611 => "111000010100001010000",
		612 => "111000010100001010000",
		613 => "111000010100001010000",
		614 => "111000010100001010000",
		615 => "111000010100001010000",
		616 => "111000010100001010000",
		617 => "111000010100001010000",
		618 => "111000010100001010000",
		619 => "111000010100001010000",
		620 => "111000010100001010000",
		621 => "111000010100001010000",
		622 => "111000010100001010000",
		623 => "111000010100001010000",
		624 => "111000010100001010000",
		625 => "111000010100001010000",
		626 => "111000010100001010000",
		627 => "111000010100001010000",
		628 => "111000010100001010000",
		629 => "111000010100001010000",
		630 => "111000010100001010000",
		631 => "111000010100001010000",
		632 => "111000010100001010000",
		633 => "111000010100001010000",
		634 => "111000010100001010000",
		635 => "111000010100001010000",
		636 => "111000010100001010000",
		637 => "111000010100001010000",
		638 => "111000010100001010000",
		639 => "111000010100001010000",
		640 => "111000010100001010000",
		641 => "111000010100001010000",
		642 => "111000010100001010000",
		643 => "111000010100001010000",
		644 => "111000010100001010000",
		645 => "111000010100001010000",
		646 => "111000010100001010000",
		647 => "111000010100001010000",
		648 => "111000010100001010000",
		649 => "111000010100001010000",
		650 => "111000010100001010000",
		651 => "111000010100001010000",
		652 => "111000010100001010000",
		653 => "111000010100001010000",
		654 => "111000010100001010000",
		655 => "111000010100001010000",
		656 => "111000010100001010000",
		657 => "111000010100001010000",
		658 => "111000010100001010000",
		659 => "111000010100001010000",
		660 => "111000010100001010000",
		661 => "111000010100001010000",
		662 => "111000010100001010000",
		663 => "111000010100001010000",
		664 => "111000010100001010000",
		665 => "111000010100001010000",
		666 => "111000010100001010000",
		667 => "111000010100001010000",
		668 => "111000010100001010000",
		669 => "111000010100001010000",
		670 => "111000010100001010000",
		671 => "111000010100001010000",
		672 => "111000010100001010000",
		673 => "111000010100001010000",
		674 => "111000010100001010000",
		675 => "111000010100001010000",
		676 => "111000010100001010000",
		677 => "111000010100001010000",
		678 => "111000010100001010000",
		679 => "111000010100001010000",
		680 => "111000010100001010000",
		681 => "111000010100001010000",
		682 => "111000010100001010000",
		683 => "111000010100001010000",
		684 => "111000010100001010000",
		685 => "111000010100001010000",
		686 => "111000010100001010000",
		687 => "111000010100001010000",
		688 => "111000010100001010000",
		689 => "111000010100001010000",
		690 => "111000010100001010000",
		691 => "111000010100001010000",
		692 => "111000010100001010000",
		693 => "111000010100001010000",
		694 => "111000010100001010000",
		695 => "111000010100001010000",
		696 => "111000010100001010000",
		697 => "111000010100001010000",
		698 => "111000010100001010000",
		699 => "111000010100001010000",
		700 => "111000010100001010000",
		701 => "111000010100001010000",
		702 => "111000010100001010000",
		703 => "111000010100001010000",
		704 => "111000010100001010000",
		705 => "111000010100001010000",
		706 => "111000010100001010000",
		707 => "111000010100001010000",
		708 => "111000010100001010000",
		709 => "111000010100001010000",
		710 => "111000010100001010000",
		711 => "111000010100001010000",
		712 => "111000010100001010000",
		713 => "111000010100001010000",
		714 => "111000010100001010000",
		715 => "111000010100001010000",
		716 => "111000010100001010000",
		717 => "111000010100001010000",
		718 => "111000010100001010000",
		719 => "111000010100001010000",
		720 => "111000010100001010000",
		721 => "111000010100001010000",
		722 => "111000010100001010000",
		723 => "111000010100001010000",
		724 => "111000010100001010000",
		725 => "111000010100001010000",
		726 => "111000010100001010000",
		727 => "111000010100001010000",
		728 => "111000010100001010000",
		729 => "111000010100001010000",
		730 => "111000010100001010000",
		731 => "111000010100001010000",
		732 => "111000010100001010000",
		733 => "111000010100001010000",
		734 => "111000010100001010000",
		735 => "111000010100001010000",
		736 => "111000010100001010000",
		737 => "111000010100001010000",
		738 => "111000010100001010000",
		739 => "111000010100001010000",
		740 => "111000010100001010000",
		741 => "111000010100001010000",
		742 => "111000010100001010000",
		743 => "111000010100001010000",
		744 => "111000010100001010000",
		745 => "111000010100001010000",
		746 => "111000010100001010000",
		747 => "111000010100001010000",
		748 => "111000010100001010000",
		749 => "111000010100001010000",
		750 => "111000010100001010000",
		751 => "111000010100001010000",
		752 => "111000010100001010000",
		753 => "111000010100001010000",
		754 => "111000010100001010000",
		755 => "111000010100001010000",
		756 => "111000010100001010000",
		757 => "111000010100001010000",
		758 => "111000010100001010000",
		759 => "111000010100001010000",
		760 => "111000010100001010000",
		761 => "111000010100001010000",
		762 => "111000010100001010000",
		763 => "111000010100001010000",
		764 => "111000010100001010000",
		765 => "111000010100001010000",
		766 => "111000010100001010000",
		767 => "111000010100001010000",
		768 => "111000010100001010000",
		769 => "111000010100001010000",
		770 => "111000010100001010000",
		771 => "111000010100001010000",
		772 => "111000010100001010000",
		773 => "111000010100001010000",
		774 => "111000010100001010000",
		775 => "111000010100001010000",
		776 => "111000010100001010000",
		777 => "111000010100001010000",
		778 => "111000010100001010000",
		779 => "111000010100001010000",
		780 => "111000010100001010000",
		781 => "111000010100001010000",
		782 => "111000010100001010000",
		783 => "111000010100001010000",
		784 => "111000010100001010000",
		785 => "111000010100001010000",
		786 => "111000010100001010000",
		787 => "111000010100001010000",
		788 => "111000010100001010000",
		789 => "111000010100001010000",
		790 => "111000010100001010000",
		791 => "111000010100001010000",
		792 => "111000010100001010000",
		793 => "111000010100001010000",
		794 => "111000010100001010000",
		795 => "111000010100001010000",
		796 => "111000010100001010000",
		797 => "111000010100001010000",
		798 => "111000010100001010000",
		799 => "111000010100001010000",
		800 => "111000010100001010000",
		801 => "111000010100001010000",
		802 => "111000010100001010000",
		803 => "111000010100001010000",
		804 => "111000010100001010000",
		805 => "111000010100001010000",
		806 => "111000010100001010000",
		807 => "111000010100001010000",
		808 => "111000010100001010000",
		809 => "111000010100001010000",
		810 => "111000010100001010000",
		811 => "111000010100001010000",
		812 => "111000010100001010000",
		813 => "111000010100001010000",
		814 => "111000010100001010000",
		815 => "111000010100001010000",
		816 => "111000010100001010000",
		817 => "111000010100001010000",
		818 => "111000010100001010000",
		819 => "111000010100001010000",
		820 => "111000010100001010000",
		821 => "111000010100001010000",
		822 => "111000010100001010000",
		823 => "111000010100001010000",
		824 => "111000010100001010000",
		825 => "111000010100001010000",
		826 => "111000010100001010000",
		827 => "111000010100001010000",
		828 => "111000010100001010000",
		829 => "111000010100001010000",
		830 => "111000010100001010000",
		831 => "111000010100001010000",
		832 => "111000010100001010000",
		833 => "111000010100001010000",
		834 => "111000010100001010000",
		835 => "111000010100001010000",
		836 => "111000010100001010000",
		837 => "111000010100001010000",
		838 => "111000010100001010000",
		839 => "111000010100001010000",
		840 => "111000010100001010000",
		841 => "111000010100001010000",
		842 => "111000010100001010000",
		843 => "111000010100001010000",
		844 => "111000010100001010000",
		845 => "111000010100001010000",
		846 => "111000010100001010000",
		847 => "111000010100001010000",
		848 => "111000010100001010000",
		849 => "111000010100001010000",
		850 => "111000010100001010000",
		851 => "111000010100001010000",
		852 => "111000010100001010000",
		853 => "111000010100001010000",
		854 => "111000010100001010000",
		855 => "111000010100001010000",
		856 => "111000010100001010000",
		857 => "111000010100001010000",
		858 => "111000010100001010000",
		859 => "111000010100001010000",
		860 => "111000010100001010000",
		861 => "111000010100001010000",
		862 => "111000010100001010000",
		863 => "111000010100001010000");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;