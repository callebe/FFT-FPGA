LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.MainPackage.all;

ENTITY TESTE IS
	PORT(Clock: IN STD_LOGIC;
		  reset: IN STD_LOGIC;
		  N: IN INTEGER RANGE 0 TO 1024;
		  SF_D : OUT STD_LOGIC_VECTOR(3 downto 0);
		  LCD_E: OUT STD_LOGIC;
		  LCD_RS: OUT STD_LOGIC;
		  LCD_RW: OUT STD_LOGIC);
END TESTE;

ARCHITECTURE Logica OF TESTE IS
	SIGNAL Even: Complex := (0,2);
	SIGNAL Odd: Complex := (0,1);
	SIGNAL DATA: INFO := ("01000001","01000110","01000001","01000110","01000001","01000110","01000001","01000110","01000001","01000110","01000001","01000110","01000001","01000110","01000111","01000001","01000110","01000001","01000110","01000001","01000110","01000001","01000110","01000001","01000110","01000001","01000110","01000001","01000110","01000111","01000111","01000111");
	
	BEGIN
	
	Display: DisplayLCD PORT MAP (Clock,reset,DATA,SF_D,LCD_E,LCD_RS,LCD_RW);
	
	
END Logica;
