library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT13 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT13;

architecture Behavioral of ROMFFT13 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 14 
	constant ROM_tb : ROM := (
		0 => "001011011100001011001",
		1 => "001011011100001011001",
		2 => "001011011100001011001",
		3 => "011011100100001010011",
		4 => "011011100100001010011",
		5 => "011011100100001010011",
		6 => "011000001110100010101",
		7 => "011000001110100010101",
		8 => "011000001110100010101",
		9 => "001001011100001010111",
		10 => "001001011100001010111",
		11 => "001001011100001010111",
		12 => "011001011101001010000",
		13 => "011001011101001010000",
		14 => "011001011101001010000",
		15 => "001000111100011110010",
		16 => "001000111100011110010",
		17 => "001000111100011110010",
		18 => "011000110100011010011",
		19 => "011000110100011010011",
		20 => "011000110100011010011",
		21 => "011000011100111010000",
		22 => "011000011100111010000",
		23 => "011000011100111010000",
		24 => "001000100100111110001",
		25 => "001000100100111110001",
		26 => "001000100100111110001",
		27 => "011001001100111110000",
		28 => "011001001100111110000",
		29 => "011001001100111110000",
		30 => "011001011100001010100",
		31 => "011001011100001010100",
		32 => "011001011100001010100",
		33 => "011000000100111010001",
		34 => "011000000100111010001",
		35 => "011000000100111010001",
		36 => "011010011100001010101",
		37 => "011010011100001010101",
		38 => "011010011100001010101",
		39 => "001000000100111110010",
		40 => "001000000100111110010",
		41 => "001000000100111110010",
		42 => "011000001111010010111",
		43 => "011000001111010010111",
		44 => "011000001111010010111",
		45 => "011000011110101011000",
		46 => "011000011110101011000",
		47 => "011000011110101011000",
		48 => "011100100100001010110",
		49 => "011100100100001010110",
		50 => "011100100100001010110",
		51 => "011011100100001010011",
		52 => "011011100100001010011",
		53 => "011011100100001010011",
		54 => "011000001110100010101",
		55 => "011000001110100010101",
		56 => "011000001110100010101",
		57 => "011010100100001010011",
		58 => "011010100100001010011",
		59 => "011010100100001010011",
		60 => "011010000100001010010",
		61 => "011010000100001010010",
		62 => "011010000100001010010",
		63 => "001000111100011110010",
		64 => "001000111100011110010",
		65 => "001000111100011110010",
		66 => "001000000100101110111",
		67 => "001000000100101110111",
		68 => "001000000100101110111",
		69 => "011001000100001110100",
		70 => "011001000100001110100",
		71 => "011001000100001110100",
		72 => "001000110100011010011",
		73 => "001000110100011010011",
		74 => "001000110100011010011",
		75 => "001000011100101110011",
		76 => "001000011100101110011",
		77 => "001000011100101110011",
		78 => "011000000101001010010",
		79 => "011000000101001010010",
		80 => "011000000101001010010",
		81 => "011000000100111010001",
		82 => "011000000100111010001",
		83 => "011000000100111010001",
		84 => "011010100100001110100",
		85 => "011010100100001110100",
		86 => "011010100100001110100",
		87 => "001001010100001010011",
		88 => "001001010100001010011",
		89 => "001001010100001010011",
		90 => "011000001111010010111",
		91 => "011000001111010010111",
		92 => "011000001111010010111",
		93 => "011000011110101011000",
		94 => "011000011110101011000",
		95 => "011000011110101011000",
		96 => "011001111101111010000",
		97 => "011001111101111010000",
		98 => "011001111101111010000",
		99 => "011001001100111010000",
		100 => "011001001100111010000",
		101 => "011001001100111010000",
		102 => "011000111101001010000",
		103 => "011000111101001010000",
		104 => "011000111101001010000",
		105 => "001001011100001010011",
		106 => "001001011100001010011",
		107 => "001001011100001010011",
		108 => "001010011100011110010",
		109 => "001010011100011110010",
		110 => "001010011100011110010",
		111 => "011000000101001010100",
		112 => "011000000101001010100",
		113 => "011000000101001010100",
		114 => "011000000101101010010",
		115 => "011000000101101010010",
		116 => "011000000101101010010",
		117 => "011100001110011110000",
		118 => "011100001110011110000",
		119 => "011100001110011110000",
		120 => "011011100100001010011",
		121 => "011011100100001010011",
		122 => "011011100100001010011",
		123 => "011001100100011110000",
		124 => "011001100100011110000",
		125 => "011001100100011110000",
		126 => "011000111101001010000",
		127 => "011000111101001010000",
		128 => "011000111101001010000",
		129 => "011001100100001010010",
		130 => "011001100100001010010",
		131 => "011001100100001010010",
		132 => "011001000100001010100",
		133 => "011001000100001010100",
		134 => "011001000100001010100",
		135 => "011010000100001110100",
		136 => "011010000100001110100",
		137 => "011010000100001110100",
		138 => "011000000101101010010",
		139 => "011000000101101010010",
		140 => "011000000101101010010",
		141 => "001000011110001111001",
		142 => "001000011110001111001",
		143 => "001000011110001111001",
		144 => "011001111101111010000",
		145 => "011001111101111010000",
		146 => "011001111101111010000",
		147 => "011001001100111010000",
		148 => "011001001100111010000",
		149 => "011001001100111010000",
		150 => "011000111101001010000",
		151 => "011000111101001010000",
		152 => "011000111101001010000",
		153 => "001001011100001010011",
		154 => "001001011100001010011",
		155 => "001001011100001010011",
		156 => "001010011100011110010",
		157 => "001010011100011110010",
		158 => "001010011100011110010",
		159 => "011000000101001010100",
		160 => "011000000101001010100",
		161 => "011000000101001010100",
		162 => "011000000101101010010",
		163 => "011000000101101010010",
		164 => "011000000101101010010",
		165 => "011100001110011110000",
		166 => "011100001110011110000",
		167 => "011100001110011110000",
		168 => "011011100100001010011",
		169 => "011011100100001010011",
		170 => "011011100100001010011",
		171 => "011001100100011110000",
		172 => "011001100100011110000",
		173 => "011001100100011110000",
		174 => "011000111101001010000",
		175 => "011000111101001010000",
		176 => "011000111101001010000",
		177 => "011001100100001010010",
		178 => "011001100100001010010",
		179 => "011001100100001010010",
		180 => "011001000100001010100",
		181 => "011001000100001010100",
		182 => "011001000100001010100",
		183 => "011010000100001110100",
		184 => "011010000100001110100",
		185 => "011010000100001110100",
		186 => "011000000101101010010",
		187 => "011000000101101010010",
		188 => "011000000101101010010",
		189 => "001000011110001111001",
		190 => "001000011110001111001",
		191 => "001000011110001111001",
		192 => "001001011100001010101",
		193 => "001001011100001010101",
		194 => "001001011100001010101",
		195 => "001010011100011110010",
		196 => "001010011100011110010",
		197 => "001010011100011110010",
		198 => "011000001101100010011",
		199 => "011000001101100010011",
		200 => "011000001101100010011",
		201 => "011000011110001010110",
		202 => "011000011110001010110",
		203 => "011000011110001010110",
		204 => "011010100100001010010",
		205 => "011010100100001010010",
		206 => "011010100100001010010",
		207 => "011001000100001010100",
		208 => "011001000100001010100",
		209 => "011001000100001010100",
		210 => "011000001101100010011",
		211 => "011000001101100010011",
		212 => "011000001101100010011",
		213 => "011100000101101010000",
		214 => "011100000101101010000",
		215 => "011100000101101010000",
		216 => "001001011100001010101",
		217 => "001001011100001010101",
		218 => "001001011100001010101",
		219 => "001010011100011110010",
		220 => "001010011100011110010",
		221 => "001010011100011110010",
		222 => "011000001101100010011",
		223 => "011000001101100010011",
		224 => "011000001101100010011",
		225 => "011000011110001010110",
		226 => "011000011110001010110",
		227 => "011000011110001010110",
		228 => "011010100100001010010",
		229 => "011010100100001010010",
		230 => "011010100100001010010",
		231 => "011001000100001010100",
		232 => "011001000100001010100",
		233 => "011001000100001010100",
		234 => "011000001101100010011",
		235 => "011000001101100010011",
		236 => "011000001101100010011",
		237 => "011100000101101010000",
		238 => "011100000101101010000",
		239 => "011100000101101010000",
		240 => "001001011100001010101",
		241 => "001001011100001010101",
		242 => "001001011100001010101",
		243 => "001010011100011110010",
		244 => "001010011100011110010",
		245 => "001010011100011110010",
		246 => "011000001101100010011",
		247 => "011000001101100010011",
		248 => "011000001101100010011",
		249 => "011000011110001010110",
		250 => "011000011110001010110",
		251 => "011000011110001010110",
		252 => "011010100100001010010",
		253 => "011010100100001010010",
		254 => "011010100100001010010",
		255 => "011001000100001010100",
		256 => "011001000100001010100",
		257 => "011001000100001010100",
		258 => "011000001101100010011",
		259 => "011000001101100010011",
		260 => "011000001101100010011",
		261 => "011100000101101010000",
		262 => "011100000101101010000",
		263 => "011100000101101010000",
		264 => "001001011100001010101",
		265 => "001001011100001010101",
		266 => "001001011100001010101",
		267 => "001010011100011110010",
		268 => "001010011100011110010",
		269 => "001010011100011110010",
		270 => "011000001101100010011",
		271 => "011000001101100010011",
		272 => "011000001101100010011",
		273 => "011000011110001010110",
		274 => "011000011110001010110",
		275 => "011000011110001010110",
		276 => "011010100100001010010",
		277 => "011010100100001010010",
		278 => "011010100100001010010",
		279 => "011001000100001010100",
		280 => "011001000100001010100",
		281 => "011001000100001010100",
		282 => "011000001101100010011",
		283 => "011000001101100010011",
		284 => "011000001101100010011",
		285 => "011100000101101010000",
		286 => "011100000101101010000",
		287 => "011100000101101010000",
		288 => "001001111100001010110",
		289 => "001001111100001010110",
		290 => "001001111100001010110",
		291 => "011000010100111010110",
		292 => "011000010100111010110",
		293 => "011000010100111010110",
		294 => "011011000100001010011",
		295 => "011011000100001010011",
		296 => "011011000100001010011",
		297 => "011000000101110011001",
		298 => "011000000101110011001",
		299 => "011000000101110011001",
		300 => "001001111100001010110",
		301 => "001001111100001010110",
		302 => "001001111100001010110",
		303 => "011000010100111010110",
		304 => "011000010100111010110",
		305 => "011000010100111010110",
		306 => "011011000100001010011",
		307 => "011011000100001010011",
		308 => "011011000100001010011",
		309 => "011000000101110011001",
		310 => "011000000101110011001",
		311 => "011000000101110011001",
		312 => "001001111100001010110",
		313 => "001001111100001010110",
		314 => "001001111100001010110",
		315 => "011000010100111010110",
		316 => "011000010100111010110",
		317 => "011000010100111010110",
		318 => "011011000100001010011",
		319 => "011011000100001010011",
		320 => "011011000100001010011",
		321 => "011000000101110011001",
		322 => "011000000101110011001",
		323 => "011000000101110011001",
		324 => "001001111100001010110",
		325 => "001001111100001010110",
		326 => "001001111100001010110",
		327 => "011000010100111010110",
		328 => "011000010100111010110",
		329 => "011000010100111010110",
		330 => "011011000100001010011",
		331 => "011011000100001010011",
		332 => "011011000100001010011",
		333 => "011000000101110011001",
		334 => "011000000101110011001",
		335 => "011000000101110011001",
		336 => "001001111100001010110",
		337 => "001001111100001010110",
		338 => "001001111100001010110",
		339 => "011000010100111010110",
		340 => "011000010100111010110",
		341 => "011000010100111010110",
		342 => "011011000100001010011",
		343 => "011011000100001010011",
		344 => "011011000100001010011",
		345 => "011000000101110011001",
		346 => "011000000101110011001",
		347 => "011000000101110011001",
		348 => "001001111100001010110",
		349 => "001001111100001010110",
		350 => "001001111100001010110",
		351 => "011000010100111010110",
		352 => "011000010100111010110",
		353 => "011000010100111010110",
		354 => "011011000100001010011",
		355 => "011011000100001010011",
		356 => "011011000100001010011",
		357 => "011000000101110011001",
		358 => "011000000101110011001",
		359 => "011000000101110011001",
		360 => "001001111100001010110",
		361 => "001001111100001010110",
		362 => "001001111100001010110",
		363 => "011000010100111010110",
		364 => "011000010100111010110",
		365 => "011000010100111010110",
		366 => "011011000100001010011",
		367 => "011011000100001010011",
		368 => "011011000100001010011",
		369 => "011000000101110011001",
		370 => "011000000101110011001",
		371 => "011000000101110011001",
		372 => "001001111100001010110",
		373 => "001001111100001010110",
		374 => "001001111100001010110",
		375 => "011000010100111010110",
		376 => "011000010100111010110",
		377 => "011000010100111010110",
		378 => "011011000100001010011",
		379 => "011011000100001010011",
		380 => "011011000100001010011",
		381 => "011000000101110011001",
		382 => "011000000101110011001",
		383 => "011000000101110011001",
		384 => "011000000101011010101",
		385 => "011000000101011010101",
		386 => "011000000101011010101",
		387 => "011000000101011010101",
		388 => "011000000101011010101",
		389 => "011000000101011010101",
		390 => "011000000101011010101",
		391 => "011000000101011010101",
		392 => "011000000101011010101",
		393 => "011000000101011010101",
		394 => "011000000101011010101",
		395 => "011000000101011010101",
		396 => "011000000101011010101",
		397 => "011000000101011010101",
		398 => "011000000101011010101",
		399 => "011000000101011010101",
		400 => "011000000101011010101",
		401 => "011000000101011010101",
		402 => "011000000101011010101",
		403 => "011000000101011010101",
		404 => "011000000101011010101",
		405 => "011000000101011010101",
		406 => "011000000101011010101",
		407 => "011000000101011010101",
		408 => "011000000101011010101",
		409 => "011000000101011010101",
		410 => "011000000101011010101",
		411 => "011000000101011010101",
		412 => "011000000101011010101",
		413 => "011000000101011010101",
		414 => "011000000101011010101",
		415 => "011000000101011010101",
		416 => "011000000101011010101",
		417 => "011000000101011010101",
		418 => "011000000101011010101",
		419 => "011000000101011010101",
		420 => "011000000101011010101",
		421 => "011000000101011010101",
		422 => "011000000101011010101",
		423 => "011000000101011010101",
		424 => "011000000101011010101",
		425 => "011000000101011010101",
		426 => "011000000101011010101",
		427 => "011000000101011010101",
		428 => "011000000101011010101",
		429 => "011000000101011010101",
		430 => "011000000101011010101",
		431 => "011000000101011010101",
		432 => "011000000101011010101",
		433 => "011000000101011010101",
		434 => "011000000101011010101",
		435 => "011000000101011010101",
		436 => "011000000101011010101",
		437 => "011000000101011010101",
		438 => "011000000101011010101",
		439 => "011000000101011010101",
		440 => "011000000101011010101",
		441 => "011000000101011010101",
		442 => "011000000101011010101",
		443 => "011000000101011010101",
		444 => "011000000101011010101",
		445 => "011000000101011010101",
		446 => "011000000101011010101",
		447 => "011000000101011010101",
		448 => "011000000101011010101",
		449 => "011000000101011010101",
		450 => "011000000101011010101",
		451 => "011000000101011010101",
		452 => "011000000101011010101",
		453 => "011000000101011010101",
		454 => "011000000101011010101",
		455 => "011000000101011010101",
		456 => "011000000101011010101",
		457 => "011000000101011010101",
		458 => "011000000101011010101",
		459 => "011000000101011010101",
		460 => "011000000101011010101",
		461 => "011000000101011010101",
		462 => "011000000101011010101",
		463 => "011000000101011010101",
		464 => "011000000101011010101",
		465 => "011000000101011010101",
		466 => "011000000101011010101",
		467 => "011000000101011010101",
		468 => "011000000101011010101",
		469 => "011000000101011010101",
		470 => "011000000101011010101",
		471 => "011000000101011010101",
		472 => "011000000101011010101",
		473 => "011000000101011010101",
		474 => "011000000101011010101",
		475 => "011000000101011010101",
		476 => "011000000101011010101",
		477 => "011000000101011010101",
		478 => "011000000101011010101",
		479 => "011000000101011010101",
		480 => "011000001101100010011",
		481 => "011000001101100010011",
		482 => "011000001101100010011",
		483 => "011000001101100010011",
		484 => "011000001101100010011",
		485 => "011000001101100010011",
		486 => "011000001101100010011",
		487 => "011000001101100010011",
		488 => "011000001101100010011",
		489 => "011000001101100010011",
		490 => "011000001101100010011",
		491 => "011000001101100010011",
		492 => "011000001101100010011",
		493 => "011000001101100010011",
		494 => "011000001101100010011",
		495 => "011000001101100010011",
		496 => "011000001101100010011",
		497 => "011000001101100010011",
		498 => "011000001101100010011",
		499 => "011000001101100010011",
		500 => "011000001101100010011",
		501 => "011000001101100010011",
		502 => "011000001101100010011",
		503 => "011000001101100010011",
		504 => "011000001101100010011",
		505 => "011000001101100010011",
		506 => "011000001101100010011",
		507 => "011000001101100010011",
		508 => "011000001101100010011",
		509 => "011000001101100010011",
		510 => "011000001101100010011",
		511 => "011000001101100010011",
		512 => "011000001101100010011",
		513 => "011000001101100010011",
		514 => "011000001101100010011",
		515 => "011000001101100010011",
		516 => "011000001101100010011",
		517 => "011000001101100010011",
		518 => "011000001101100010011",
		519 => "011000001101100010011",
		520 => "011000001101100010011",
		521 => "011000001101100010011",
		522 => "011000001101100010011",
		523 => "011000001101100010011",
		524 => "011000001101100010011",
		525 => "011000001101100010011",
		526 => "011000001101100010011",
		527 => "011000001101100010011",
		528 => "011000001101100010011",
		529 => "011000001101100010011",
		530 => "011000001101100010011",
		531 => "011000001101100010011",
		532 => "011000001101100010011",
		533 => "011000001101100010011",
		534 => "011000001101100010011",
		535 => "011000001101100010011",
		536 => "011000001101100010011",
		537 => "011000001101100010011",
		538 => "011000001101100010011",
		539 => "011000001101100010011",
		540 => "011000001101100010011",
		541 => "011000001101100010011",
		542 => "011000001101100010011",
		543 => "011000001101100010011",
		544 => "011000001101100010011",
		545 => "011000001101100010011",
		546 => "011000001101100010011",
		547 => "011000001101100010011",
		548 => "011000001101100010011",
		549 => "011000001101100010011",
		550 => "011000001101100010011",
		551 => "011000001101100010011",
		552 => "011000001101100010011",
		553 => "011000001101100010011",
		554 => "011000001101100010011",
		555 => "011000001101100010011",
		556 => "011000001101100010011",
		557 => "011000001101100010011",
		558 => "011000001101100010011",
		559 => "011000001101100010011",
		560 => "011000001101100010011",
		561 => "011000001101100010011",
		562 => "011000001101100010011",
		563 => "011000001101100010011",
		564 => "011000001101100010011",
		565 => "011000001101100010011",
		566 => "011000001101100010011",
		567 => "011000001101100010011",
		568 => "011000001101100010011",
		569 => "011000001101100010011",
		570 => "011000001101100010011",
		571 => "011000001101100010011",
		572 => "011000001101100010011",
		573 => "011000001101100010011",
		574 => "011000001101100010011",
		575 => "011000001101100010011",
		576 => "011011000100001110011",
		577 => "011011000100001110011",
		578 => "011011000100001110011",
		579 => "011011000100001110011",
		580 => "011011000100001110011",
		581 => "011011000100001110011",
		582 => "011011000100001110011",
		583 => "011011000100001110011",
		584 => "011011000100001110011",
		585 => "011011000100001110011",
		586 => "011011000100001110011",
		587 => "011011000100001110011",
		588 => "011011000100001110011",
		589 => "011011000100001110011",
		590 => "011011000100001110011",
		591 => "011011000100001110011",
		592 => "011011000100001110011",
		593 => "011011000100001110011",
		594 => "011011000100001110011",
		595 => "011011000100001110011",
		596 => "011011000100001110011",
		597 => "011011000100001110011",
		598 => "011011000100001110011",
		599 => "011011000100001110011",
		600 => "011011000100001110011",
		601 => "011011000100001110011",
		602 => "011011000100001110011",
		603 => "011011000100001110011",
		604 => "011011000100001110011",
		605 => "011011000100001110011",
		606 => "011011000100001110011",
		607 => "011011000100001110011",
		608 => "011011000100001110011",
		609 => "011011000100001110011",
		610 => "011011000100001110011",
		611 => "011011000100001110011",
		612 => "011011000100001110011",
		613 => "011011000100001110011",
		614 => "011011000100001110011",
		615 => "011011000100001110011",
		616 => "011011000100001110011",
		617 => "011011000100001110011",
		618 => "011011000100001110011",
		619 => "011011000100001110011",
		620 => "011011000100001110011",
		621 => "011011000100001110011",
		622 => "011011000100001110011",
		623 => "011011000100001110011",
		624 => "011011000100001110011",
		625 => "011011000100001110011",
		626 => "011011000100001110011",
		627 => "011011000100001110011",
		628 => "011011000100001110011",
		629 => "011011000100001110011",
		630 => "011011000100001110011",
		631 => "011011000100001110011",
		632 => "011011000100001110011",
		633 => "011011000100001110011",
		634 => "011011000100001110011",
		635 => "011011000100001110011",
		636 => "011011000100001110011",
		637 => "011011000100001110011",
		638 => "011011000100001110011",
		639 => "011011000100001110011",
		640 => "011011000100001110011",
		641 => "011011000100001110011",
		642 => "011011000100001110011",
		643 => "011011000100001110011",
		644 => "011011000100001110011",
		645 => "011011000100001110011",
		646 => "011011000100001110011",
		647 => "011011000100001110011",
		648 => "011011000100001110011",
		649 => "011011000100001110011",
		650 => "011011000100001110011",
		651 => "011011000100001110011",
		652 => "011011000100001110011",
		653 => "011011000100001110011",
		654 => "011011000100001110011",
		655 => "011011000100001110011",
		656 => "011011000100001110011",
		657 => "011011000100001110011",
		658 => "011011000100001110011",
		659 => "011011000100001110011",
		660 => "011011000100001110011",
		661 => "011011000100001110011",
		662 => "011011000100001110011",
		663 => "011011000100001110011",
		664 => "011011000100001110011",
		665 => "011011000100001110011",
		666 => "011011000100001110011",
		667 => "011011000100001110011",
		668 => "011011000100001110011",
		669 => "011011000100001110011",
		670 => "011011000100001110011",
		671 => "011011000100001110011",
		672 => "011000101100100010101",
		673 => "011000101100100010101",
		674 => "011000101100100010101",
		675 => "011000101100100010101",
		676 => "011000101100100010101",
		677 => "011000101100100010101",
		678 => "011000101100100010101",
		679 => "011000101100100010101",
		680 => "011000101100100010101",
		681 => "011000101100100010101",
		682 => "011000101100100010101",
		683 => "011000101100100010101",
		684 => "011000101100100010101",
		685 => "011000101100100010101",
		686 => "011000101100100010101",
		687 => "011000101100100010101",
		688 => "011000101100100010101",
		689 => "011000101100100010101",
		690 => "011000101100100010101",
		691 => "011000101100100010101",
		692 => "011000101100100010101",
		693 => "011000101100100010101",
		694 => "011000101100100010101",
		695 => "011000101100100010101",
		696 => "011000101100100010101",
		697 => "011000101100100010101",
		698 => "011000101100100010101",
		699 => "011000101100100010101",
		700 => "011000101100100010101",
		701 => "011000101100100010101",
		702 => "011000101100100010101",
		703 => "011000101100100010101",
		704 => "011000101100100010101",
		705 => "011000101100100010101",
		706 => "011000101100100010101",
		707 => "011000101100100010101",
		708 => "011000101100100010101",
		709 => "011000101100100010101",
		710 => "011000101100100010101",
		711 => "011000101100100010101",
		712 => "011000101100100010101",
		713 => "011000101100100010101",
		714 => "011000101100100010101",
		715 => "011000101100100010101",
		716 => "011000101100100010101",
		717 => "011000101100100010101",
		718 => "011000101100100010101",
		719 => "011000101100100010101",
		720 => "011000101100100010101",
		721 => "011000101100100010101",
		722 => "011000101100100010101",
		723 => "011000101100100010101",
		724 => "011000101100100010101",
		725 => "011000101100100010101",
		726 => "011000101100100010101",
		727 => "011000101100100010101",
		728 => "011000101100100010101",
		729 => "011000101100100010101",
		730 => "011000101100100010101",
		731 => "011000101100100010101",
		732 => "011000101100100010101",
		733 => "011000101100100010101",
		734 => "011000101100100010101",
		735 => "011000101100100010101",
		736 => "011000101100100010101",
		737 => "011000101100100010101",
		738 => "011000101100100010101",
		739 => "011000101100100010101",
		740 => "011000101100100010101",
		741 => "011000101100100010101",
		742 => "011000101100100010101",
		743 => "011000101100100010101",
		744 => "011000101100100010101",
		745 => "011000101100100010101",
		746 => "011000101100100010101",
		747 => "011000101100100010101",
		748 => "011000101100100010101",
		749 => "011000101100100010101",
		750 => "011000101100100010101",
		751 => "011000101100100010101",
		752 => "011000101100100010101",
		753 => "011000101100100010101",
		754 => "011000101100100010101",
		755 => "011000101100100010101",
		756 => "011000101100100010101",
		757 => "011000101100100010101",
		758 => "011000101100100010101",
		759 => "011000101100100010101",
		760 => "011000101100100010101",
		761 => "011000101100100010101",
		762 => "011000101100100010101",
		763 => "011000101100100010101",
		764 => "011000101100100010101",
		765 => "011000101100100010101",
		766 => "011000101100100010101",
		767 => "011000101100100010101",
		768 => "011000101100100110010",
		769 => "011000101100100110010",
		770 => "011000101100100110010",
		771 => "011000101100100110010",
		772 => "011000101100100110010",
		773 => "011000101100100110010",
		774 => "011000101100100110010",
		775 => "011000101100100110010",
		776 => "011000101100100110010",
		777 => "011000101100100110010",
		778 => "011000101100100110010",
		779 => "011000101100100110010",
		780 => "011000101100100110010",
		781 => "011000101100100110010",
		782 => "011000101100100110010",
		783 => "011000101100100110010",
		784 => "011000101100100110010",
		785 => "011000101100100110010",
		786 => "011000101100100110010",
		787 => "011000101100100110010",
		788 => "011000101100100110010",
		789 => "011000101100100110010",
		790 => "011000101100100110010",
		791 => "011000101100100110010",
		792 => "011000101100100110010",
		793 => "011000101100100110010",
		794 => "011000101100100110010",
		795 => "011000101100100110010",
		796 => "011000101100100110010",
		797 => "011000101100100110010",
		798 => "011000101100100110010",
		799 => "011000101100100110010",
		800 => "011000101100100110010",
		801 => "011000101100100110010",
		802 => "011000101100100110010",
		803 => "011000101100100110010",
		804 => "011000101100100110010",
		805 => "011000101100100110010",
		806 => "011000101100100110010",
		807 => "011000101100100110010",
		808 => "011000101100100110010",
		809 => "011000101100100110010",
		810 => "011000101100100110010",
		811 => "011000101100100110010",
		812 => "011000101100100110010",
		813 => "011000101100100110010",
		814 => "011000101100100110010",
		815 => "011000101100100110010",
		816 => "011000101100100110010",
		817 => "011000101100100110010",
		818 => "011000101100100110010",
		819 => "011000101100100110010",
		820 => "011000101100100110010",
		821 => "011000101100100110010",
		822 => "011000101100100110010",
		823 => "011000101100100110010",
		824 => "011000101100100110010",
		825 => "011000101100100110010",
		826 => "011000101100100110010",
		827 => "011000101100100110010",
		828 => "011000101100100110010",
		829 => "011000101100100110010",
		830 => "011000101100100110010",
		831 => "011000101100100110010",
		832 => "011000101100100110010",
		833 => "011000101100100110010",
		834 => "011000101100100110010",
		835 => "011000101100100110010",
		836 => "011000101100100110010",
		837 => "011000101100100110010",
		838 => "011000101100100110010",
		839 => "011000101100100110010",
		840 => "011000101100100110010",
		841 => "011000101100100110010",
		842 => "011000101100100110010",
		843 => "011000101100100110010",
		844 => "011000101100100110010",
		845 => "011000101100100110010",
		846 => "011000101100100110010",
		847 => "011000101100100110010",
		848 => "011000101100100110010",
		849 => "011000101100100110010",
		850 => "011000101100100110010",
		851 => "011000101100100110010",
		852 => "011000101100100110010",
		853 => "011000101100100110010",
		854 => "011000101100100110010",
		855 => "011000101100100110010",
		856 => "011000101100100110010",
		857 => "011000101100100110010",
		858 => "011000101100100110010",
		859 => "011000101100100110010",
		860 => "011000101100100110010",
		861 => "011000101100100110010",
		862 => "011000101100100110010",
		863 => "011000101100100110010");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;