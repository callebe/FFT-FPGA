library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT1024p_7 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT1024p_7;

architecture Behavioral of ROMFFT1024p_7 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 8 
	constant ROM_tb : ROM := (
		0 => "001010100101111110000",
		1 => "001010100101111110000",
		2 => "001010100101111110000",
		3 => "001010111100001011001",
		4 => "001010111100001011001",
		5 => "001010111100001011001",
		6 => "011011100100001010110",
		7 => "011011100100001010110",
		8 => "011011100100001010110",
		9 => "001001111100001010110",
		10 => "001001111100001010110",
		11 => "001001111100001010110",
		12 => "011011111100001010101",
		13 => "011011111100001010101",
		14 => "011011111100001010101",
		15 => "001010111100001010101",
		16 => "001010111100001010101",
		17 => "001010111100001010101",
		18 => "011010100100101110000",
		19 => "011010100100101110000",
		20 => "011010100100101110000",
		21 => "011000000100111110001",
		22 => "011000000100111110001",
		23 => "011000000100111110001",
		24 => "011000110100001010101",
		25 => "011000110100001010101",
		26 => "011000110100001010101",
		27 => "011000101100101010001",
		28 => "011000101100101010001",
		29 => "011000101100101010001",
		30 => "011000111100111010000",
		31 => "011000111100111010000",
		32 => "011000111100111010000",
		33 => "001000111100001010011",
		34 => "001000111100001010011",
		35 => "001000111100001010011",
		36 => "011000000100111010000",
		37 => "011000000100111010000",
		38 => "011000000100111010000",
		39 => "001000111100011110011",
		40 => "001000111100011110011",
		41 => "001000111100011110011",
		42 => "011000101100111110001",
		43 => "011000101100111110001",
		44 => "011000101100111110001",
		45 => "001000111100001010011",
		46 => "001000111100001010011",
		47 => "001000111100001010011",
		48 => "001001011100111010000",
		49 => "001001011100111010000",
		50 => "001001011100111010000",
		51 => "011000101100111010001",
		52 => "011000101100111010001",
		53 => "011000101100111010001",
		54 => "011000111100011110011",
		55 => "011000111100011110011",
		56 => "011000111100011110011",
		57 => "011000001100110010110",
		58 => "011000001100110010110",
		59 => "011000001100110010110",
		60 => "011001111100001010100",
		61 => "011001111100001010100",
		62 => "011001111100001010100",
		63 => "011000000101001010010",
		64 => "011000000101001010010",
		65 => "011000000101001010010",
		66 => "011000001101100010011",
		67 => "011000001101100010011",
		68 => "011000001101100010011",
		69 => "011001100100001110001",
		70 => "011001100100001110001",
		71 => "011001100100001110001",
		72 => "011001000100001110001",
		73 => "011001000100001110001",
		74 => "011001000100001110001",
		75 => "011000000101011010100",
		76 => "011000000101011010100",
		77 => "011000000101011010100",
		78 => "011001011100001010101",
		79 => "011001011100001010101",
		80 => "011001011100001010101",
		81 => "011000010100111010110",
		82 => "011000010100111010110",
		83 => "011000010100111010110",
		84 => "011000000101101010011",
		85 => "011000000101101010011",
		86 => "011000000101101010011",
		87 => "001011011100001010111",
		88 => "001011011100001010111",
		89 => "001011011100001010111",
		90 => "011100100100001110100",
		91 => "011100100100001110100",
		92 => "011100100100001110100",
		93 => "011100100111001010000",
		94 => "011100100111001010000",
		95 => "011100100111001010000",
		96 => "011011100101001110000",
		97 => "011011100101001110000",
		98 => "011011100101001110000",
		99 => "001010011100001010111",
		100 => "001010011100001010111",
		101 => "001010011100001010111",
		102 => "001001111100001010101",
		103 => "001001111100001010101",
		104 => "001001111100001010101",
		105 => "011000110100001010010",
		106 => "011000110100001010010",
		107 => "011000110100001010010",
		108 => "001011011100001010011",
		109 => "001011011100001010011",
		110 => "001011011100001010011",
		111 => "001000100100111110000",
		112 => "001000100100111110000",
		113 => "001000100100111110000",
		114 => "001000111100011110011",
		115 => "001000111100011110011",
		116 => "001000111100011110011",
		117 => "011000011100111010000",
		118 => "011000011100111010000",
		119 => "011000011100111010000",
		120 => "011000001100101010101",
		121 => "011000001100101010101",
		122 => "011000001100101010101",
		123 => "011001111100001010011",
		124 => "011001111100001010011",
		125 => "011001111100001010011",
		126 => "011000000101011010010",
		127 => "011000000101011010010",
		128 => "011000000101011010010",
		129 => "011001100100001110010",
		130 => "011001100100001110010",
		131 => "011001100100001110010",
		132 => "011010100100001110100",
		133 => "011010100100001110100",
		134 => "011010100100001110100",
		135 => "001010111100001010101",
		136 => "001010111100001010101",
		137 => "001010111100001010101",
		138 => "011011011101111010000",
		139 => "011011011101111010000",
		140 => "011011011101111010000",
		141 => "001000011101101011011",
		142 => "001000011101101011011",
		143 => "001000011101101011011",
		144 => "001000011101111010100",
		145 => "001000011101111010100",
		146 => "001000011101111010100",
		147 => "011011100100001010100",
		148 => "011011100100001010100",
		149 => "011011100100001010100",
		150 => "011010100100001010011",
		151 => "011010100100001010011",
		152 => "011010100100001010011",
		153 => "001000111100001110010",
		154 => "001000111100001110010",
		155 => "001000111100001110010",
		156 => "011001100100001010110",
		157 => "011001100100001010110",
		158 => "011001100100001010110",
		159 => "001000010100011010011",
		160 => "001000010100011010011",
		161 => "001000010100011010011",
		162 => "001000100100111010001",
		163 => "001000100100111010001",
		164 => "001000100100111010001",
		165 => "011001000100001110100",
		166 => "011001000100001110100",
		167 => "011001000100001110100",
		168 => "001000100100111110001",
		169 => "001000100100111110001",
		170 => "001000100100111110001",
		171 => "011001100100001110011",
		172 => "011001100100001110011",
		173 => "011001100100001110011",
		174 => "011000000101011010010",
		175 => "011000000101011010010",
		176 => "011000000101011010010",
		177 => "011000000100111010010",
		178 => "011000000100111010010",
		179 => "011000000100111010010",
		180 => "011010100100001110100",
		181 => "011010100100001110100",
		182 => "011010100100001110100",
		183 => "011010100100001010101",
		184 => "011010100100001010101",
		185 => "011010100100001010101",
		186 => "011011100100001010110",
		187 => "011011100100001010110",
		188 => "011011100100001010110",
		189 => "011101100101101010000",
		190 => "011101100101101010000",
		191 => "011101100101101010000",
		192 => "001010011100001010111",
		193 => "001010011100001010111",
		194 => "001010011100001010111",
		195 => "011010100100001010010",
		196 => "011010100100001010010",
		197 => "011010100100001010010",
		198 => "001001011100001010100",
		199 => "001001011100001010100",
		200 => "001001011100001010100",
		201 => "011000011100111010000",
		202 => "011000011100111010000",
		203 => "011000011100111010000",
		204 => "001001111100011110010",
		205 => "001001111100011110010",
		206 => "001001111100011110010",
		207 => "001000110100001010011",
		208 => "001000110100001010011",
		209 => "001000110100001010011",
		210 => "011000000101011010010",
		211 => "011000000101011010010",
		212 => "011000000101011010010",
		213 => "011000000110111010101",
		214 => "011000000110111010101",
		215 => "011000000110111010101",
		216 => "001000011101101010011",
		217 => "001000011101101010011",
		218 => "001000011101101010011",
		219 => "011010100100001010010",
		220 => "011010100100001010010",
		221 => "011010100100001010010",
		222 => "011010000100001010010",
		223 => "011010000100001010010",
		224 => "011010000100001010010",
		225 => "011001000100001110100",
		226 => "011001000100001110100",
		227 => "011001000100001110100",
		228 => "011001000100001010011",
		229 => "011001000100001010011",
		230 => "011001000100001010011",
		231 => "011000101100100110100",
		232 => "011000101100100110100",
		233 => "011000101100100110100",
		234 => "001001011101011010000",
		235 => "001001011101011010000",
		236 => "001001011101011010000",
		237 => "001000011110101010111",
		238 => "001000011110101010111",
		239 => "001000011110101010111",
		240 => "001010011100001010111",
		241 => "001010011100001010111",
		242 => "001010011100001010111",
		243 => "011010100100001010010",
		244 => "011010100100001010010",
		245 => "011010100100001010010",
		246 => "001001011100001010100",
		247 => "001001011100001010100",
		248 => "001001011100001010100",
		249 => "011000011100111010000",
		250 => "011000011100111010000",
		251 => "011000011100111010000",
		252 => "001001111100011110010",
		253 => "001001111100011110010",
		254 => "001001111100011110010",
		255 => "001000110100001010011",
		256 => "001000110100001010011",
		257 => "001000110100001010011",
		258 => "011000000101011010010",
		259 => "011000000101011010010",
		260 => "011000000101011010010",
		261 => "011000000110111010101",
		262 => "011000000110111010101",
		263 => "011000000110111010101",
		264 => "001000011101101010011",
		265 => "001000011101101010011",
		266 => "001000011101101010011",
		267 => "011010100100001010010",
		268 => "011010100100001010010",
		269 => "011010100100001010010",
		270 => "011010000100001010010",
		271 => "011010000100001010010",
		272 => "011010000100001010010",
		273 => "011001000100001110100",
		274 => "011001000100001110100",
		275 => "011001000100001110100",
		276 => "011001000100001010011",
		277 => "011001000100001010011",
		278 => "011001000100001010011",
		279 => "011000101100100110100",
		280 => "011000101100100110100",
		281 => "011000101100100110100",
		282 => "001001011101011010000",
		283 => "001001011101011010000",
		284 => "001001011101011010000",
		285 => "001000011110101010111",
		286 => "001000011110101010111",
		287 => "001000011110101010111",
		288 => "001001111100001010101",
		289 => "001001111100001010101",
		290 => "001001111100001010101",
		291 => "011001011100111010000",
		292 => "011001011100111010000",
		293 => "011001011100111010000",
		294 => "011000001101110010011",
		295 => "011000001101110010011",
		296 => "011000001101110010011",
		297 => "011000000110011010100",
		298 => "011000000110011010100",
		299 => "011000000110011010100",
		300 => "001000011101011010010",
		301 => "001000011101011010010",
		302 => "001000011101011010010",
		303 => "011001100100001010010",
		304 => "011001100100001010010",
		305 => "011001100100001010010",
		306 => "011000001101110010011",
		307 => "011000001101110010011",
		308 => "011000001101110010011",
		309 => "001010011110011010000",
		310 => "001010011110011010000",
		311 => "001010011110011010000",
		312 => "001001111100001010101",
		313 => "001001111100001010101",
		314 => "001001111100001010101",
		315 => "011001011100111010000",
		316 => "011001011100111010000",
		317 => "011001011100111010000",
		318 => "011000001101110010011",
		319 => "011000001101110010011",
		320 => "011000001101110010011",
		321 => "011000000110011010100",
		322 => "011000000110011010100",
		323 => "011000000110011010100",
		324 => "001000011101011010010",
		325 => "001000011101011010010",
		326 => "001000011101011010010",
		327 => "011001100100001010010",
		328 => "011001100100001010010",
		329 => "011001100100001010010",
		330 => "011000001101110010011",
		331 => "011000001101110010011",
		332 => "011000001101110010011",
		333 => "001010011110011010000",
		334 => "001010011110011010000",
		335 => "001010011110011010000",
		336 => "001001111100001010101",
		337 => "001001111100001010101",
		338 => "001001111100001010101",
		339 => "011001011100111010000",
		340 => "011001011100111010000",
		341 => "011001011100111010000",
		342 => "011000001101110010011",
		343 => "011000001101110010011",
		344 => "011000001101110010011",
		345 => "011000000110011010100",
		346 => "011000000110011010100",
		347 => "011000000110011010100",
		348 => "001000011101011010010",
		349 => "001000011101011010010",
		350 => "001000011101011010010",
		351 => "011001100100001010010",
		352 => "011001100100001010010",
		353 => "011001100100001010010",
		354 => "011000001101110010011",
		355 => "011000001101110010011",
		356 => "011000001101110010011",
		357 => "001010011110011010000",
		358 => "001010011110011010000",
		359 => "001010011110011010000",
		360 => "001001111100001010101",
		361 => "001001111100001010101",
		362 => "001001111100001010101",
		363 => "011001011100111010000",
		364 => "011001011100111010000",
		365 => "011001011100111010000",
		366 => "011000001101110010011",
		367 => "011000001101110010011",
		368 => "011000001101110010011",
		369 => "011000000110011010100",
		370 => "011000000110011010100",
		371 => "011000000110011010100",
		372 => "001000011101011010010",
		373 => "001000011101011010010",
		374 => "001000011101011010010",
		375 => "011001100100001010010",
		376 => "011001100100001010010",
		377 => "011001100100001010010",
		378 => "011000001101110010011",
		379 => "011000001101110010011",
		380 => "011000001101110010011",
		381 => "001010011110011010000",
		382 => "001010011110011010000",
		383 => "001010011110011010000",
		384 => "001000111100011110011",
		385 => "001000111100011110011",
		386 => "001000111100011110011",
		387 => "011011100100001110011",
		388 => "011011100100001110011",
		389 => "011011100100001110011",
		390 => "001000100100111010001",
		391 => "001000100100111010001",
		392 => "001000100100111010001",
		393 => "011000000101111010011",
		394 => "011000000101111010011",
		395 => "011000000101111010011",
		396 => "001000111100011110011",
		397 => "001000111100011110011",
		398 => "001000111100011110011",
		399 => "011011100100001110011",
		400 => "011011100100001110011",
		401 => "011011100100001110011",
		402 => "001000100100111010001",
		403 => "001000100100111010001",
		404 => "001000100100111010001",
		405 => "011000000101111010011",
		406 => "011000000101111010011",
		407 => "011000000101111010011",
		408 => "001000111100011110011",
		409 => "001000111100011110011",
		410 => "001000111100011110011",
		411 => "011011100100001110011",
		412 => "011011100100001110011",
		413 => "011011100100001110011",
		414 => "001000100100111010001",
		415 => "001000100100111010001",
		416 => "001000100100111010001",
		417 => "011000000101111010011",
		418 => "011000000101111010011",
		419 => "011000000101111010011",
		420 => "001000111100011110011",
		421 => "001000111100011110011",
		422 => "001000111100011110011",
		423 => "011011100100001110011",
		424 => "011011100100001110011",
		425 => "011011100100001110011",
		426 => "001000100100111010001",
		427 => "001000100100111010001",
		428 => "001000100100111010001",
		429 => "011000000101111010011",
		430 => "011000000101111010011",
		431 => "011000000101111010011",
		432 => "001000111100011110011",
		433 => "001000111100011110011",
		434 => "001000111100011110011",
		435 => "011011100100001110011",
		436 => "011011100100001110011",
		437 => "011011100100001110011",
		438 => "001000100100111010001",
		439 => "001000100100111010001",
		440 => "001000100100111010001",
		441 => "011000000101111010011",
		442 => "011000000101111010011",
		443 => "011000000101111010011",
		444 => "001000111100011110011",
		445 => "001000111100011110011",
		446 => "001000111100011110011",
		447 => "011011100100001110011",
		448 => "011011100100001110011",
		449 => "011011100100001110011",
		450 => "001000100100111010001",
		451 => "001000100100111010001",
		452 => "001000100100111010001",
		453 => "011000000101111010011",
		454 => "011000000101111010011",
		455 => "011000000101111010011",
		456 => "001000111100011110011",
		457 => "001000111100011110011",
		458 => "001000111100011110011",
		459 => "011011100100001110011",
		460 => "011011100100001110011",
		461 => "011011100100001110011",
		462 => "001000100100111010001",
		463 => "001000100100111010001",
		464 => "001000100100111010001",
		465 => "011000000101111010011",
		466 => "011000000101111010011",
		467 => "011000000101111010011",
		468 => "001000111100011110011",
		469 => "001000111100011110011",
		470 => "001000111100011110011",
		471 => "011011100100001110011",
		472 => "011011100100001110011",
		473 => "011011100100001110011",
		474 => "001000100100111010001",
		475 => "001000100100111010001",
		476 => "001000100100111010001",
		477 => "011000000101111010011",
		478 => "011000000101111010011",
		479 => "011000000101111010011",
		480 => "011010100100001010100",
		481 => "011010100100001010100",
		482 => "011010100100001010100",
		483 => "011010100100001010100",
		484 => "011010100100001010100",
		485 => "011010100100001010100",
		486 => "011010100100001010100",
		487 => "011010100100001010100",
		488 => "011010100100001010100",
		489 => "011010100100001010100",
		490 => "011010100100001010100",
		491 => "011010100100001010100",
		492 => "011010100100001010100",
		493 => "011010100100001010100",
		494 => "011010100100001010100",
		495 => "011010100100001010100",
		496 => "011010100100001010100",
		497 => "011010100100001010100",
		498 => "011010100100001010100",
		499 => "011010100100001010100",
		500 => "011010100100001010100",
		501 => "011010100100001010100",
		502 => "011010100100001010100",
		503 => "011010100100001010100",
		504 => "011010100100001010100",
		505 => "011010100100001010100",
		506 => "011010100100001010100",
		507 => "011010100100001010100",
		508 => "011010100100001010100",
		509 => "011010100100001010100",
		510 => "011010100100001010100",
		511 => "011010100100001010100",
		512 => "011010100100001010100",
		513 => "011010100100001010100",
		514 => "011010100100001010100",
		515 => "011010100100001010100",
		516 => "011010100100001010100",
		517 => "011010100100001010100",
		518 => "011010100100001010100",
		519 => "011010100100001010100",
		520 => "011010100100001010100",
		521 => "011010100100001010100",
		522 => "011010100100001010100",
		523 => "011010100100001010100",
		524 => "011010100100001010100",
		525 => "011010100100001010100",
		526 => "011010100100001010100",
		527 => "011010100100001010100",
		528 => "011010100100001010100",
		529 => "011010100100001010100",
		530 => "011010100100001010100",
		531 => "011010100100001010100",
		532 => "011010100100001010100",
		533 => "011010100100001010100",
		534 => "011010100100001010100",
		535 => "011010100100001010100",
		536 => "011010100100001010100",
		537 => "011010100100001010100",
		538 => "011010100100001010100",
		539 => "011010100100001010100",
		540 => "011010100100001010100",
		541 => "011010100100001010100",
		542 => "011010100100001010100",
		543 => "011010100100001010100",
		544 => "011010100100001010100",
		545 => "011010100100001010100",
		546 => "011010100100001010100",
		547 => "011010100100001010100",
		548 => "011010100100001010100",
		549 => "011010100100001010100",
		550 => "011010100100001010100",
		551 => "011010100100001010100",
		552 => "011010100100001010100",
		553 => "011010100100001010100",
		554 => "011010100100001010100",
		555 => "011010100100001010100",
		556 => "011010100100001010100",
		557 => "011010100100001010100",
		558 => "011010100100001010100",
		559 => "011010100100001010100",
		560 => "011010100100001010100",
		561 => "011010100100001010100",
		562 => "011010100100001010100",
		563 => "011010100100001010100",
		564 => "011010100100001010100",
		565 => "011010100100001010100",
		566 => "011010100100001010100",
		567 => "011010100100001010100",
		568 => "011010100100001010100",
		569 => "011010100100001010100",
		570 => "011010100100001010100",
		571 => "011010100100001010100",
		572 => "011010100100001010100",
		573 => "011010100100001010100",
		574 => "011010100100001010100",
		575 => "011010100100001010100",
		576 => "001000111100111010000",
		577 => "001000111100111010000",
		578 => "001000111100111010000",
		579 => "001000111100111010000",
		580 => "001000111100111010000",
		581 => "001000111100111010000",
		582 => "001000111100111010000",
		583 => "001000111100111010000",
		584 => "001000111100111010000",
		585 => "001000111100111010000",
		586 => "001000111100111010000",
		587 => "001000111100111010000",
		588 => "001000111100111010000",
		589 => "001000111100111010000",
		590 => "001000111100111010000",
		591 => "001000111100111010000",
		592 => "001000111100111010000",
		593 => "001000111100111010000",
		594 => "001000111100111010000",
		595 => "001000111100111010000",
		596 => "001000111100111010000",
		597 => "001000111100111010000",
		598 => "001000111100111010000",
		599 => "001000111100111010000",
		600 => "001000111100111010000",
		601 => "001000111100111010000",
		602 => "001000111100111010000",
		603 => "001000111100111010000",
		604 => "001000111100111010000",
		605 => "001000111100111010000",
		606 => "001000111100111010000",
		607 => "001000111100111010000",
		608 => "001000111100111010000",
		609 => "001000111100111010000",
		610 => "001000111100111010000",
		611 => "001000111100111010000",
		612 => "001000111100111010000",
		613 => "001000111100111010000",
		614 => "001000111100111010000",
		615 => "001000111100111010000",
		616 => "001000111100111010000",
		617 => "001000111100111010000",
		618 => "001000111100111010000",
		619 => "001000111100111010000",
		620 => "001000111100111010000",
		621 => "001000111100111010000",
		622 => "001000111100111010000",
		623 => "001000111100111010000",
		624 => "001000111100111010000",
		625 => "001000111100111010000",
		626 => "001000111100111010000",
		627 => "001000111100111010000",
		628 => "001000111100111010000",
		629 => "001000111100111010000",
		630 => "001000111100111010000",
		631 => "001000111100111010000",
		632 => "001000111100111010000",
		633 => "001000111100111010000",
		634 => "001000111100111010000",
		635 => "001000111100111010000",
		636 => "001000111100111010000",
		637 => "001000111100111010000",
		638 => "001000111100111010000",
		639 => "001000111100111010000",
		640 => "001000111100111010000",
		641 => "001000111100111010000",
		642 => "001000111100111010000",
		643 => "001000111100111010000",
		644 => "001000111100111010000",
		645 => "001000111100111010000",
		646 => "001000111100111010000",
		647 => "001000111100111010000",
		648 => "001000111100111010000",
		649 => "001000111100111010000",
		650 => "001000111100111010000",
		651 => "001000111100111010000",
		652 => "001000111100111010000",
		653 => "001000111100111010000",
		654 => "001000111100111010000",
		655 => "001000111100111010000",
		656 => "001000111100111010000",
		657 => "001000111100111010000",
		658 => "001000111100111010000",
		659 => "001000111100111010000",
		660 => "001000111100111010000",
		661 => "001000111100111010000",
		662 => "001000111100111010000",
		663 => "001000111100111010000",
		664 => "001000111100111010000",
		665 => "001000111100111010000",
		666 => "001000111100111010000",
		667 => "001000111100111010000",
		668 => "001000111100111010000",
		669 => "001000111100111010000",
		670 => "001000111100111010000",
		671 => "001000111100111010000",
		672 => "011000101100100010101",
		673 => "011000101100100010101",
		674 => "011000101100100010101",
		675 => "011000101100100010101",
		676 => "011000101100100010101",
		677 => "011000101100100010101",
		678 => "011000101100100010101",
		679 => "011000101100100010101",
		680 => "011000101100100010101",
		681 => "011000101100100010101",
		682 => "011000101100100010101",
		683 => "011000101100100010101",
		684 => "011000101100100010101",
		685 => "011000101100100010101",
		686 => "011000101100100010101",
		687 => "011000101100100010101",
		688 => "011000101100100010101",
		689 => "011000101100100010101",
		690 => "011000101100100010101",
		691 => "011000101100100010101",
		692 => "011000101100100010101",
		693 => "011000101100100010101",
		694 => "011000101100100010101",
		695 => "011000101100100010101",
		696 => "011000101100100010101",
		697 => "011000101100100010101",
		698 => "011000101100100010101",
		699 => "011000101100100010101",
		700 => "011000101100100010101",
		701 => "011000101100100010101",
		702 => "011000101100100010101",
		703 => "011000101100100010101",
		704 => "011000101100100010101",
		705 => "011000101100100010101",
		706 => "011000101100100010101",
		707 => "011000101100100010101",
		708 => "011000101100100010101",
		709 => "011000101100100010101",
		710 => "011000101100100010101",
		711 => "011000101100100010101",
		712 => "011000101100100010101",
		713 => "011000101100100010101",
		714 => "011000101100100010101",
		715 => "011000101100100010101",
		716 => "011000101100100010101",
		717 => "011000101100100010101",
		718 => "011000101100100010101",
		719 => "011000101100100010101",
		720 => "011000101100100010101",
		721 => "011000101100100010101",
		722 => "011000101100100010101",
		723 => "011000101100100010101",
		724 => "011000101100100010101",
		725 => "011000101100100010101",
		726 => "011000101100100010101",
		727 => "011000101100100010101",
		728 => "011000101100100010101",
		729 => "011000101100100010101",
		730 => "011000101100100010101",
		731 => "011000101100100010101",
		732 => "011000101100100010101",
		733 => "011000101100100010101",
		734 => "011000101100100010101",
		735 => "011000101100100010101",
		736 => "011000101100100010101",
		737 => "011000101100100010101",
		738 => "011000101100100010101",
		739 => "011000101100100010101",
		740 => "011000101100100010101",
		741 => "011000101100100010101",
		742 => "011000101100100010101",
		743 => "011000101100100010101",
		744 => "011000101100100010101",
		745 => "011000101100100010101",
		746 => "011000101100100010101",
		747 => "011000101100100010101",
		748 => "011000101100100010101",
		749 => "011000101100100010101",
		750 => "011000101100100010101",
		751 => "011000101100100010101",
		752 => "011000101100100010101",
		753 => "011000101100100010101",
		754 => "011000101100100010101",
		755 => "011000101100100010101",
		756 => "011000101100100010101",
		757 => "011000101100100010101",
		758 => "011000101100100010101",
		759 => "011000101100100010101",
		760 => "011000101100100010101",
		761 => "011000101100100010101",
		762 => "011000101100100010101",
		763 => "011000101100100010101",
		764 => "011000101100100010101",
		765 => "011000101100100010101",
		766 => "011000101100100010101",
		767 => "011000101100100010101",
		768 => "011000101100100110010",
		769 => "011000101100100110010",
		770 => "011000101100100110010",
		771 => "011000101100100110010",
		772 => "011000101100100110010",
		773 => "011000101100100110010",
		774 => "011000101100100110010",
		775 => "011000101100100110010",
		776 => "011000101100100110010",
		777 => "011000101100100110010",
		778 => "011000101100100110010",
		779 => "011000101100100110010",
		780 => "011000101100100110010",
		781 => "011000101100100110010",
		782 => "011000101100100110010",
		783 => "011000101100100110010",
		784 => "011000101100100110010",
		785 => "011000101100100110010",
		786 => "011000101100100110010",
		787 => "011000101100100110010",
		788 => "011000101100100110010",
		789 => "011000101100100110010",
		790 => "011000101100100110010",
		791 => "011000101100100110010",
		792 => "011000101100100110010",
		793 => "011000101100100110010",
		794 => "011000101100100110010",
		795 => "011000101100100110010",
		796 => "011000101100100110010",
		797 => "011000101100100110010",
		798 => "011000101100100110010",
		799 => "011000101100100110010",
		800 => "011000101100100110010",
		801 => "011000101100100110010",
		802 => "011000101100100110010",
		803 => "011000101100100110010",
		804 => "011000101100100110010",
		805 => "011000101100100110010",
		806 => "011000101100100110010",
		807 => "011000101100100110010",
		808 => "011000101100100110010",
		809 => "011000101100100110010",
		810 => "011000101100100110010",
		811 => "011000101100100110010",
		812 => "011000101100100110010",
		813 => "011000101100100110010",
		814 => "011000101100100110010",
		815 => "011000101100100110010",
		816 => "011000101100100110010",
		817 => "011000101100100110010",
		818 => "011000101100100110010",
		819 => "011000101100100110010",
		820 => "011000101100100110010",
		821 => "011000101100100110010",
		822 => "011000101100100110010",
		823 => "011000101100100110010",
		824 => "011000101100100110010",
		825 => "011000101100100110010",
		826 => "011000101100100110010",
		827 => "011000101100100110010",
		828 => "011000101100100110010",
		829 => "011000101100100110010",
		830 => "011000101100100110010",
		831 => "011000101100100110010",
		832 => "011000101100100110010",
		833 => "011000101100100110010",
		834 => "011000101100100110010",
		835 => "011000101100100110010",
		836 => "011000101100100110010",
		837 => "011000101100100110010",
		838 => "011000101100100110010",
		839 => "011000101100100110010",
		840 => "011000101100100110010",
		841 => "011000101100100110010",
		842 => "011000101100100110010",
		843 => "011000101100100110010",
		844 => "011000101100100110010",
		845 => "011000101100100110010",
		846 => "011000101100100110010",
		847 => "011000101100100110010",
		848 => "011000101100100110010",
		849 => "011000101100100110010",
		850 => "011000101100100110010",
		851 => "011000101100100110010",
		852 => "011000101100100110010",
		853 => "011000101100100110010",
		854 => "011000101100100110010",
		855 => "011000101100100110010",
		856 => "011000101100100110010",
		857 => "011000101100100110010",
		858 => "011000101100100110010",
		859 => "011000101100100110010",
		860 => "011000101100100110010",
		861 => "011000101100100110010",
		862 => "011000101100100110010",
		863 => "011000101100100110010");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;