library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT14 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT14;

architecture Behavioral of ROMFFT14 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 15 
	constant ROM_tb : ROM := (
		0 => "011011100101001110000",
		1 => "011011100101001110000",
		2 => "011011100101001110000",
		3 => "001010011100001010111",
		4 => "001010011100001010111",
		5 => "001010011100001010111",
		6 => "001001111100001010101",
		7 => "001001111100001010101",
		8 => "001001111100001010101",
		9 => "011000110100001010010",
		10 => "011000110100001010010",
		11 => "011000110100001010010",
		12 => "001011011100001010011",
		13 => "001011011100001010011",
		14 => "001011011100001010011",
		15 => "001000100100111110000",
		16 => "001000100100111110000",
		17 => "001000100100111110000",
		18 => "001000111100011110011",
		19 => "001000111100011110011",
		20 => "001000111100011110011",
		21 => "011000011100111010000",
		22 => "011000011100111010000",
		23 => "011000011100111010000",
		24 => "011000001100101010101",
		25 => "011000001100101010101",
		26 => "011000001100101010101",
		27 => "011001111100001010011",
		28 => "011001111100001010011",
		29 => "011001111100001010011",
		30 => "011000000101011010010",
		31 => "011000000101011010010",
		32 => "011000000101011010010",
		33 => "011001100100001110010",
		34 => "011001100100001110010",
		35 => "011001100100001110010",
		36 => "011010100100001110100",
		37 => "011010100100001110100",
		38 => "011010100100001110100",
		39 => "001010111100001010101",
		40 => "001010111100001010101",
		41 => "001010111100001010101",
		42 => "011011011101111010000",
		43 => "011011011101111010000",
		44 => "011011011101111010000",
		45 => "001000011101101011011",
		46 => "001000011101101011011",
		47 => "001000011101101011011",
		48 => "001000011101111010100",
		49 => "001000011101111010100",
		50 => "001000011101111010100",
		51 => "011011100100001010100",
		52 => "011011100100001010100",
		53 => "011011100100001010100",
		54 => "011010100100001010011",
		55 => "011010100100001010011",
		56 => "011010100100001010011",
		57 => "001000111100001110010",
		58 => "001000111100001110010",
		59 => "001000111100001110010",
		60 => "011001100100001010110",
		61 => "011001100100001010110",
		62 => "011001100100001010110",
		63 => "001000010100011010011",
		64 => "001000010100011010011",
		65 => "001000010100011010011",
		66 => "001000100100111010001",
		67 => "001000100100111010001",
		68 => "001000100100111010001",
		69 => "011001000100001110100",
		70 => "011001000100001110100",
		71 => "011001000100001110100",
		72 => "001000100100111110001",
		73 => "001000100100111110001",
		74 => "001000100100111110001",
		75 => "011001100100001110011",
		76 => "011001100100001110011",
		77 => "011001100100001110011",
		78 => "011000000101011010010",
		79 => "011000000101011010010",
		80 => "011000000101011010010",
		81 => "011000000100111010010",
		82 => "011000000100111010010",
		83 => "011000000100111010010",
		84 => "011010100100001110100",
		85 => "011010100100001110100",
		86 => "011010100100001110100",
		87 => "011010100100001010101",
		88 => "011010100100001010101",
		89 => "011010100100001010101",
		90 => "011011100100001010110",
		91 => "011011100100001010110",
		92 => "011011100100001010110",
		93 => "011101100101101010000",
		94 => "011101100101101010000",
		95 => "011101100101101010000",
		96 => "001010011100001010111",
		97 => "001010011100001010111",
		98 => "001010011100001010111",
		99 => "011010100100001010010",
		100 => "011010100100001010010",
		101 => "011010100100001010010",
		102 => "001001011100001010100",
		103 => "001001011100001010100",
		104 => "001001011100001010100",
		105 => "011000011100111010000",
		106 => "011000011100111010000",
		107 => "011000011100111010000",
		108 => "001001111100011110010",
		109 => "001001111100011110010",
		110 => "001001111100011110010",
		111 => "001000110100001010011",
		112 => "001000110100001010011",
		113 => "001000110100001010011",
		114 => "011000000101011010010",
		115 => "011000000101011010010",
		116 => "011000000101011010010",
		117 => "011000000110111010101",
		118 => "011000000110111010101",
		119 => "011000000110111010101",
		120 => "001000011101101010011",
		121 => "001000011101101010011",
		122 => "001000011101101010011",
		123 => "011010100100001010010",
		124 => "011010100100001010010",
		125 => "011010100100001010010",
		126 => "011010000100001010010",
		127 => "011010000100001010010",
		128 => "011010000100001010010",
		129 => "011001000100001110100",
		130 => "011001000100001110100",
		131 => "011001000100001110100",
		132 => "011001000100001010011",
		133 => "011001000100001010011",
		134 => "011001000100001010011",
		135 => "011000101100100110100",
		136 => "011000101100100110100",
		137 => "011000101100100110100",
		138 => "001001011101011010000",
		139 => "001001011101011010000",
		140 => "001001011101011010000",
		141 => "001000011110101010111",
		142 => "001000011110101010111",
		143 => "001000011110101010111",
		144 => "001010011100001010111",
		145 => "001010011100001010111",
		146 => "001010011100001010111",
		147 => "011010100100001010010",
		148 => "011010100100001010010",
		149 => "011010100100001010010",
		150 => "001001011100001010100",
		151 => "001001011100001010100",
		152 => "001001011100001010100",
		153 => "011000011100111010000",
		154 => "011000011100111010000",
		155 => "011000011100111010000",
		156 => "001001111100011110010",
		157 => "001001111100011110010",
		158 => "001001111100011110010",
		159 => "001000110100001010011",
		160 => "001000110100001010011",
		161 => "001000110100001010011",
		162 => "011000000101011010010",
		163 => "011000000101011010010",
		164 => "011000000101011010010",
		165 => "011000000110111010101",
		166 => "011000000110111010101",
		167 => "011000000110111010101",
		168 => "001000011101101010011",
		169 => "001000011101101010011",
		170 => "001000011101101010011",
		171 => "011010100100001010010",
		172 => "011010100100001010010",
		173 => "011010100100001010010",
		174 => "011010000100001010010",
		175 => "011010000100001010010",
		176 => "011010000100001010010",
		177 => "011001000100001110100",
		178 => "011001000100001110100",
		179 => "011001000100001110100",
		180 => "011001000100001010011",
		181 => "011001000100001010011",
		182 => "011001000100001010011",
		183 => "011000101100100110100",
		184 => "011000101100100110100",
		185 => "011000101100100110100",
		186 => "001001011101011010000",
		187 => "001001011101011010000",
		188 => "001001011101011010000",
		189 => "001000011110101010111",
		190 => "001000011110101010111",
		191 => "001000011110101010111",
		192 => "001001111100001010101",
		193 => "001001111100001010101",
		194 => "001001111100001010101",
		195 => "011001011100111010000",
		196 => "011001011100111010000",
		197 => "011001011100111010000",
		198 => "011000001101110010011",
		199 => "011000001101110010011",
		200 => "011000001101110010011",
		201 => "011000000110011010100",
		202 => "011000000110011010100",
		203 => "011000000110011010100",
		204 => "001000011101011010010",
		205 => "001000011101011010010",
		206 => "001000011101011010010",
		207 => "011001100100001010010",
		208 => "011001100100001010010",
		209 => "011001100100001010010",
		210 => "011000001101110010011",
		211 => "011000001101110010011",
		212 => "011000001101110010011",
		213 => "001010011110011010000",
		214 => "001010011110011010000",
		215 => "001010011110011010000",
		216 => "001001111100001010101",
		217 => "001001111100001010101",
		218 => "001001111100001010101",
		219 => "011001011100111010000",
		220 => "011001011100111010000",
		221 => "011001011100111010000",
		222 => "011000001101110010011",
		223 => "011000001101110010011",
		224 => "011000001101110010011",
		225 => "011000000110011010100",
		226 => "011000000110011010100",
		227 => "011000000110011010100",
		228 => "001000011101011010010",
		229 => "001000011101011010010",
		230 => "001000011101011010010",
		231 => "011001100100001010010",
		232 => "011001100100001010010",
		233 => "011001100100001010010",
		234 => "011000001101110010011",
		235 => "011000001101110010011",
		236 => "011000001101110010011",
		237 => "001010011110011010000",
		238 => "001010011110011010000",
		239 => "001010011110011010000",
		240 => "001001111100001010101",
		241 => "001001111100001010101",
		242 => "001001111100001010101",
		243 => "011001011100111010000",
		244 => "011001011100111010000",
		245 => "011001011100111010000",
		246 => "011000001101110010011",
		247 => "011000001101110010011",
		248 => "011000001101110010011",
		249 => "011000000110011010100",
		250 => "011000000110011010100",
		251 => "011000000110011010100",
		252 => "001000011101011010010",
		253 => "001000011101011010010",
		254 => "001000011101011010010",
		255 => "011001100100001010010",
		256 => "011001100100001010010",
		257 => "011001100100001010010",
		258 => "011000001101110010011",
		259 => "011000001101110010011",
		260 => "011000001101110010011",
		261 => "001010011110011010000",
		262 => "001010011110011010000",
		263 => "001010011110011010000",
		264 => "001001111100001010101",
		265 => "001001111100001010101",
		266 => "001001111100001010101",
		267 => "011001011100111010000",
		268 => "011001011100111010000",
		269 => "011001011100111010000",
		270 => "011000001101110010011",
		271 => "011000001101110010011",
		272 => "011000001101110010011",
		273 => "011000000110011010100",
		274 => "011000000110011010100",
		275 => "011000000110011010100",
		276 => "001000011101011010010",
		277 => "001000011101011010010",
		278 => "001000011101011010010",
		279 => "011001100100001010010",
		280 => "011001100100001010010",
		281 => "011001100100001010010",
		282 => "011000001101110010011",
		283 => "011000001101110010011",
		284 => "011000001101110010011",
		285 => "001010011110011010000",
		286 => "001010011110011010000",
		287 => "001010011110011010000",
		288 => "001000111100011110011",
		289 => "001000111100011110011",
		290 => "001000111100011110011",
		291 => "011011100100001110011",
		292 => "011011100100001110011",
		293 => "011011100100001110011",
		294 => "001000100100111010001",
		295 => "001000100100111010001",
		296 => "001000100100111010001",
		297 => "011000000101111010011",
		298 => "011000000101111010011",
		299 => "011000000101111010011",
		300 => "001000111100011110011",
		301 => "001000111100011110011",
		302 => "001000111100011110011",
		303 => "011011100100001110011",
		304 => "011011100100001110011",
		305 => "011011100100001110011",
		306 => "001000100100111010001",
		307 => "001000100100111010001",
		308 => "001000100100111010001",
		309 => "011000000101111010011",
		310 => "011000000101111010011",
		311 => "011000000101111010011",
		312 => "001000111100011110011",
		313 => "001000111100011110011",
		314 => "001000111100011110011",
		315 => "011011100100001110011",
		316 => "011011100100001110011",
		317 => "011011100100001110011",
		318 => "001000100100111010001",
		319 => "001000100100111010001",
		320 => "001000100100111010001",
		321 => "011000000101111010011",
		322 => "011000000101111010011",
		323 => "011000000101111010011",
		324 => "001000111100011110011",
		325 => "001000111100011110011",
		326 => "001000111100011110011",
		327 => "011011100100001110011",
		328 => "011011100100001110011",
		329 => "011011100100001110011",
		330 => "001000100100111010001",
		331 => "001000100100111010001",
		332 => "001000100100111010001",
		333 => "011000000101111010011",
		334 => "011000000101111010011",
		335 => "011000000101111010011",
		336 => "001000111100011110011",
		337 => "001000111100011110011",
		338 => "001000111100011110011",
		339 => "011011100100001110011",
		340 => "011011100100001110011",
		341 => "011011100100001110011",
		342 => "001000100100111010001",
		343 => "001000100100111010001",
		344 => "001000100100111010001",
		345 => "011000000101111010011",
		346 => "011000000101111010011",
		347 => "011000000101111010011",
		348 => "001000111100011110011",
		349 => "001000111100011110011",
		350 => "001000111100011110011",
		351 => "011011100100001110011",
		352 => "011011100100001110011",
		353 => "011011100100001110011",
		354 => "001000100100111010001",
		355 => "001000100100111010001",
		356 => "001000100100111010001",
		357 => "011000000101111010011",
		358 => "011000000101111010011",
		359 => "011000000101111010011",
		360 => "001000111100011110011",
		361 => "001000111100011110011",
		362 => "001000111100011110011",
		363 => "011011100100001110011",
		364 => "011011100100001110011",
		365 => "011011100100001110011",
		366 => "001000100100111010001",
		367 => "001000100100111010001",
		368 => "001000100100111010001",
		369 => "011000000101111010011",
		370 => "011000000101111010011",
		371 => "011000000101111010011",
		372 => "001000111100011110011",
		373 => "001000111100011110011",
		374 => "001000111100011110011",
		375 => "011011100100001110011",
		376 => "011011100100001110011",
		377 => "011011100100001110011",
		378 => "001000100100111010001",
		379 => "001000100100111010001",
		380 => "001000100100111010001",
		381 => "011000000101111010011",
		382 => "011000000101111010011",
		383 => "011000000101111010011",
		384 => "011010100100001010100",
		385 => "011010100100001010100",
		386 => "011010100100001010100",
		387 => "011010100100001010100",
		388 => "011010100100001010100",
		389 => "011010100100001010100",
		390 => "011010100100001010100",
		391 => "011010100100001010100",
		392 => "011010100100001010100",
		393 => "011010100100001010100",
		394 => "011010100100001010100",
		395 => "011010100100001010100",
		396 => "011010100100001010100",
		397 => "011010100100001010100",
		398 => "011010100100001010100",
		399 => "011010100100001010100",
		400 => "011010100100001010100",
		401 => "011010100100001010100",
		402 => "011010100100001010100",
		403 => "011010100100001010100",
		404 => "011010100100001010100",
		405 => "011010100100001010100",
		406 => "011010100100001010100",
		407 => "011010100100001010100",
		408 => "011010100100001010100",
		409 => "011010100100001010100",
		410 => "011010100100001010100",
		411 => "011010100100001010100",
		412 => "011010100100001010100",
		413 => "011010100100001010100",
		414 => "011010100100001010100",
		415 => "011010100100001010100",
		416 => "011010100100001010100",
		417 => "011010100100001010100",
		418 => "011010100100001010100",
		419 => "011010100100001010100",
		420 => "011010100100001010100",
		421 => "011010100100001010100",
		422 => "011010100100001010100",
		423 => "011010100100001010100",
		424 => "011010100100001010100",
		425 => "011010100100001010100",
		426 => "011010100100001010100",
		427 => "011010100100001010100",
		428 => "011010100100001010100",
		429 => "011010100100001010100",
		430 => "011010100100001010100",
		431 => "011010100100001010100",
		432 => "011010100100001010100",
		433 => "011010100100001010100",
		434 => "011010100100001010100",
		435 => "011010100100001010100",
		436 => "011010100100001010100",
		437 => "011010100100001010100",
		438 => "011010100100001010100",
		439 => "011010100100001010100",
		440 => "011010100100001010100",
		441 => "011010100100001010100",
		442 => "011010100100001010100",
		443 => "011010100100001010100",
		444 => "011010100100001010100",
		445 => "011010100100001010100",
		446 => "011010100100001010100",
		447 => "011010100100001010100",
		448 => "011010100100001010100",
		449 => "011010100100001010100",
		450 => "011010100100001010100",
		451 => "011010100100001010100",
		452 => "011010100100001010100",
		453 => "011010100100001010100",
		454 => "011010100100001010100",
		455 => "011010100100001010100",
		456 => "011010100100001010100",
		457 => "011010100100001010100",
		458 => "011010100100001010100",
		459 => "011010100100001010100",
		460 => "011010100100001010100",
		461 => "011010100100001010100",
		462 => "011010100100001010100",
		463 => "011010100100001010100",
		464 => "011010100100001010100",
		465 => "011010100100001010100",
		466 => "011010100100001010100",
		467 => "011010100100001010100",
		468 => "011010100100001010100",
		469 => "011010100100001010100",
		470 => "011010100100001010100",
		471 => "011010100100001010100",
		472 => "011010100100001010100",
		473 => "011010100100001010100",
		474 => "011010100100001010100",
		475 => "011010100100001010100",
		476 => "011010100100001010100",
		477 => "011010100100001010100",
		478 => "011010100100001010100",
		479 => "011010100100001010100",
		480 => "001000111100111010000",
		481 => "001000111100111010000",
		482 => "001000111100111010000",
		483 => "001000111100111010000",
		484 => "001000111100111010000",
		485 => "001000111100111010000",
		486 => "001000111100111010000",
		487 => "001000111100111010000",
		488 => "001000111100111010000",
		489 => "001000111100111010000",
		490 => "001000111100111010000",
		491 => "001000111100111010000",
		492 => "001000111100111010000",
		493 => "001000111100111010000",
		494 => "001000111100111010000",
		495 => "001000111100111010000",
		496 => "001000111100111010000",
		497 => "001000111100111010000",
		498 => "001000111100111010000",
		499 => "001000111100111010000",
		500 => "001000111100111010000",
		501 => "001000111100111010000",
		502 => "001000111100111010000",
		503 => "001000111100111010000",
		504 => "001000111100111010000",
		505 => "001000111100111010000",
		506 => "001000111100111010000",
		507 => "001000111100111010000",
		508 => "001000111100111010000",
		509 => "001000111100111010000",
		510 => "001000111100111010000",
		511 => "001000111100111010000",
		512 => "001000111100111010000",
		513 => "001000111100111010000",
		514 => "001000111100111010000",
		515 => "001000111100111010000",
		516 => "001000111100111010000",
		517 => "001000111100111010000",
		518 => "001000111100111010000",
		519 => "001000111100111010000",
		520 => "001000111100111010000",
		521 => "001000111100111010000",
		522 => "001000111100111010000",
		523 => "001000111100111010000",
		524 => "001000111100111010000",
		525 => "001000111100111010000",
		526 => "001000111100111010000",
		527 => "001000111100111010000",
		528 => "001000111100111010000",
		529 => "001000111100111010000",
		530 => "001000111100111010000",
		531 => "001000111100111010000",
		532 => "001000111100111010000",
		533 => "001000111100111010000",
		534 => "001000111100111010000",
		535 => "001000111100111010000",
		536 => "001000111100111010000",
		537 => "001000111100111010000",
		538 => "001000111100111010000",
		539 => "001000111100111010000",
		540 => "001000111100111010000",
		541 => "001000111100111010000",
		542 => "001000111100111010000",
		543 => "001000111100111010000",
		544 => "001000111100111010000",
		545 => "001000111100111010000",
		546 => "001000111100111010000",
		547 => "001000111100111010000",
		548 => "001000111100111010000",
		549 => "001000111100111010000",
		550 => "001000111100111010000",
		551 => "001000111100111010000",
		552 => "001000111100111010000",
		553 => "001000111100111010000",
		554 => "001000111100111010000",
		555 => "001000111100111010000",
		556 => "001000111100111010000",
		557 => "001000111100111010000",
		558 => "001000111100111010000",
		559 => "001000111100111010000",
		560 => "001000111100111010000",
		561 => "001000111100111010000",
		562 => "001000111100111010000",
		563 => "001000111100111010000",
		564 => "001000111100111010000",
		565 => "001000111100111010000",
		566 => "001000111100111010000",
		567 => "001000111100111010000",
		568 => "001000111100111010000",
		569 => "001000111100111010000",
		570 => "001000111100111010000",
		571 => "001000111100111010000",
		572 => "001000111100111010000",
		573 => "001000111100111010000",
		574 => "001000111100111010000",
		575 => "001000111100111010000",
		576 => "011000101100100010101",
		577 => "011000101100100010101",
		578 => "011000101100100010101",
		579 => "011000101100100010101",
		580 => "011000101100100010101",
		581 => "011000101100100010101",
		582 => "011000101100100010101",
		583 => "011000101100100010101",
		584 => "011000101100100010101",
		585 => "011000101100100010101",
		586 => "011000101100100010101",
		587 => "011000101100100010101",
		588 => "011000101100100010101",
		589 => "011000101100100010101",
		590 => "011000101100100010101",
		591 => "011000101100100010101",
		592 => "011000101100100010101",
		593 => "011000101100100010101",
		594 => "011000101100100010101",
		595 => "011000101100100010101",
		596 => "011000101100100010101",
		597 => "011000101100100010101",
		598 => "011000101100100010101",
		599 => "011000101100100010101",
		600 => "011000101100100010101",
		601 => "011000101100100010101",
		602 => "011000101100100010101",
		603 => "011000101100100010101",
		604 => "011000101100100010101",
		605 => "011000101100100010101",
		606 => "011000101100100010101",
		607 => "011000101100100010101",
		608 => "011000101100100010101",
		609 => "011000101100100010101",
		610 => "011000101100100010101",
		611 => "011000101100100010101",
		612 => "011000101100100010101",
		613 => "011000101100100010101",
		614 => "011000101100100010101",
		615 => "011000101100100010101",
		616 => "011000101100100010101",
		617 => "011000101100100010101",
		618 => "011000101100100010101",
		619 => "011000101100100010101",
		620 => "011000101100100010101",
		621 => "011000101100100010101",
		622 => "011000101100100010101",
		623 => "011000101100100010101",
		624 => "011000101100100010101",
		625 => "011000101100100010101",
		626 => "011000101100100010101",
		627 => "011000101100100010101",
		628 => "011000101100100010101",
		629 => "011000101100100010101",
		630 => "011000101100100010101",
		631 => "011000101100100010101",
		632 => "011000101100100010101",
		633 => "011000101100100010101",
		634 => "011000101100100010101",
		635 => "011000101100100010101",
		636 => "011000101100100010101",
		637 => "011000101100100010101",
		638 => "011000101100100010101",
		639 => "011000101100100010101",
		640 => "011000101100100010101",
		641 => "011000101100100010101",
		642 => "011000101100100010101",
		643 => "011000101100100010101",
		644 => "011000101100100010101",
		645 => "011000101100100010101",
		646 => "011000101100100010101",
		647 => "011000101100100010101",
		648 => "011000101100100010101",
		649 => "011000101100100010101",
		650 => "011000101100100010101",
		651 => "011000101100100010101",
		652 => "011000101100100010101",
		653 => "011000101100100010101",
		654 => "011000101100100010101",
		655 => "011000101100100010101",
		656 => "011000101100100010101",
		657 => "011000101100100010101",
		658 => "011000101100100010101",
		659 => "011000101100100010101",
		660 => "011000101100100010101",
		661 => "011000101100100010101",
		662 => "011000101100100010101",
		663 => "011000101100100010101",
		664 => "011000101100100010101",
		665 => "011000101100100010101",
		666 => "011000101100100010101",
		667 => "011000101100100010101",
		668 => "011000101100100010101",
		669 => "011000101100100010101",
		670 => "011000101100100010101",
		671 => "011000101100100010101",
		672 => "011000101100100110010",
		673 => "011000101100100110010",
		674 => "011000101100100110010",
		675 => "011000101100100110010",
		676 => "011000101100100110010",
		677 => "011000101100100110010",
		678 => "011000101100100110010",
		679 => "011000101100100110010",
		680 => "011000101100100110010",
		681 => "011000101100100110010",
		682 => "011000101100100110010",
		683 => "011000101100100110010",
		684 => "011000101100100110010",
		685 => "011000101100100110010",
		686 => "011000101100100110010",
		687 => "011000101100100110010",
		688 => "011000101100100110010",
		689 => "011000101100100110010",
		690 => "011000101100100110010",
		691 => "011000101100100110010",
		692 => "011000101100100110010",
		693 => "011000101100100110010",
		694 => "011000101100100110010",
		695 => "011000101100100110010",
		696 => "011000101100100110010",
		697 => "011000101100100110010",
		698 => "011000101100100110010",
		699 => "011000101100100110010",
		700 => "011000101100100110010",
		701 => "011000101100100110010",
		702 => "011000101100100110010",
		703 => "011000101100100110010",
		704 => "011000101100100110010",
		705 => "011000101100100110010",
		706 => "011000101100100110010",
		707 => "011000101100100110010",
		708 => "011000101100100110010",
		709 => "011000101100100110010",
		710 => "011000101100100110010",
		711 => "011000101100100110010",
		712 => "011000101100100110010",
		713 => "011000101100100110010",
		714 => "011000101100100110010",
		715 => "011000101100100110010",
		716 => "011000101100100110010",
		717 => "011000101100100110010",
		718 => "011000101100100110010",
		719 => "011000101100100110010",
		720 => "011000101100100110010",
		721 => "011000101100100110010",
		722 => "011000101100100110010",
		723 => "011000101100100110010",
		724 => "011000101100100110010",
		725 => "011000101100100110010",
		726 => "011000101100100110010",
		727 => "011000101100100110010",
		728 => "011000101100100110010",
		729 => "011000101100100110010",
		730 => "011000101100100110010",
		731 => "011000101100100110010",
		732 => "011000101100100110010",
		733 => "011000101100100110010",
		734 => "011000101100100110010",
		735 => "011000101100100110010",
		736 => "011000101100100110010",
		737 => "011000101100100110010",
		738 => "011000101100100110010",
		739 => "011000101100100110010",
		740 => "011000101100100110010",
		741 => "011000101100100110010",
		742 => "011000101100100110010",
		743 => "011000101100100110010",
		744 => "011000101100100110010",
		745 => "011000101100100110010",
		746 => "011000101100100110010",
		747 => "011000101100100110010",
		748 => "011000101100100110010",
		749 => "011000101100100110010",
		750 => "011000101100100110010",
		751 => "011000101100100110010",
		752 => "011000101100100110010",
		753 => "011000101100100110010",
		754 => "011000101100100110010",
		755 => "011000101100100110010",
		756 => "011000101100100110010",
		757 => "011000101100100110010",
		758 => "011000101100100110010",
		759 => "011000101100100110010",
		760 => "011000101100100110010",
		761 => "011000101100100110010",
		762 => "011000101100100110010",
		763 => "011000101100100110010",
		764 => "011000101100100110010",
		765 => "011000101100100110010",
		766 => "011000101100100110010",
		767 => "011000101100100110010",
		768 => "111000010100001010000",
		769 => "111000010100001010000",
		770 => "111000010100001010000",
		771 => "111000010100001010000",
		772 => "111000010100001010000",
		773 => "111000010100001010000",
		774 => "111000010100001010000",
		775 => "111000010100001010000",
		776 => "111000010100001010000",
		777 => "111000010100001010000",
		778 => "111000010100001010000",
		779 => "111000010100001010000",
		780 => "111000010100001010000",
		781 => "111000010100001010000",
		782 => "111000010100001010000",
		783 => "111000010100001010000",
		784 => "111000010100001010000",
		785 => "111000010100001010000",
		786 => "111000010100001010000",
		787 => "111000010100001010000",
		788 => "111000010100001010000",
		789 => "111000010100001010000",
		790 => "111000010100001010000",
		791 => "111000010100001010000",
		792 => "111000010100001010000",
		793 => "111000010100001010000",
		794 => "111000010100001010000",
		795 => "111000010100001010000",
		796 => "111000010100001010000",
		797 => "111000010100001010000",
		798 => "111000010100001010000",
		799 => "111000010100001010000",
		800 => "111000010100001010000",
		801 => "111000010100001010000",
		802 => "111000010100001010000",
		803 => "111000010100001010000",
		804 => "111000010100001010000",
		805 => "111000010100001010000",
		806 => "111000010100001010000",
		807 => "111000010100001010000",
		808 => "111000010100001010000",
		809 => "111000010100001010000",
		810 => "111000010100001010000",
		811 => "111000010100001010000",
		812 => "111000010100001010000",
		813 => "111000010100001010000",
		814 => "111000010100001010000",
		815 => "111000010100001010000",
		816 => "111000010100001010000",
		817 => "111000010100001010000",
		818 => "111000010100001010000",
		819 => "111000010100001010000",
		820 => "111000010100001010000",
		821 => "111000010100001010000",
		822 => "111000010100001010000",
		823 => "111000010100001010000",
		824 => "111000010100001010000",
		825 => "111000010100001010000",
		826 => "111000010100001010000",
		827 => "111000010100001010000",
		828 => "111000010100001010000",
		829 => "111000010100001010000",
		830 => "111000010100001010000",
		831 => "111000010100001010000",
		832 => "111000010100001010000",
		833 => "111000010100001010000",
		834 => "111000010100001010000",
		835 => "111000010100001010000",
		836 => "111000010100001010000",
		837 => "111000010100001010000",
		838 => "111000010100001010000",
		839 => "111000010100001010000",
		840 => "111000010100001010000",
		841 => "111000010100001010000",
		842 => "111000010100001010000",
		843 => "111000010100001010000",
		844 => "111000010100001010000",
		845 => "111000010100001010000",
		846 => "111000010100001010000",
		847 => "111000010100001010000",
		848 => "111000010100001010000",
		849 => "111000010100001010000",
		850 => "111000010100001010000",
		851 => "111000010100001010000",
		852 => "111000010100001010000",
		853 => "111000010100001010000",
		854 => "111000010100001010000",
		855 => "111000010100001010000",
		856 => "111000010100001010000",
		857 => "111000010100001010000",
		858 => "111000010100001010000",
		859 => "111000010100001010000",
		860 => "111000010100001010000",
		861 => "111000010100001010000",
		862 => "111000010100001010000",
		863 => "111000010100001010000");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;