library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT5 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT5;

architecture Behavioral of ROMFFT5 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 6 
	constant ROM_tb : ROM := (
		0 => "001101111110111010000",
		1 => "001101111110111010000",
		2 => "001101111110111010000",
		3 => "001010000110001110000",
		4 => "001010000110001110000",
		5 => "001010000110001110000",
		6 => "011011011100001010101",
		7 => "011011011100001010101",
		8 => "011011011100001010101",
		9 => "001010011100001010101",
		10 => "001010011100001010101",
		11 => "001010011100001010101",
		12 => "011010000100001010001",
		13 => "011010000100001010001",
		14 => "011010000100001010001",
		15 => "011000000100111110001",
		16 => "011000000100111110001",
		17 => "011000000100111110001",
		18 => "011000101100101010011",
		19 => "011000101100101010011",
		20 => "011000101100101010011",
		21 => "011000000100111010000",
		22 => "011000000100111010000",
		23 => "011000000100111010000",
		24 => "001001011100111010000",
		25 => "001001011100111010000",
		26 => "001001011100111010000",
		27 => "011000011100111010000",
		28 => "011000011100111010000",
		29 => "011000011100111010000",
		30 => "011000000100111010001",
		31 => "011000000100111010001",
		32 => "011000000100111010001",
		33 => "001011011100001010011",
		34 => "001011011100001010011",
		35 => "001011011100001010011",
		36 => "001000011100011110101",
		37 => "001000011100011110101",
		38 => "001000011100011110101",
		39 => "011000000101101010010",
		40 => "011000000101101010010",
		41 => "011000000101101010010",
		42 => "011000101100101010011",
		43 => "011000101100101010011",
		44 => "011000101100101010011",
		45 => "011000000110011011000",
		46 => "011000000110011011000",
		47 => "011000000110011011000",
		48 => "011101100100001111011",
		49 => "011101100100001111011",
		50 => "011101100100001111011",
		51 => "011000000110010011100",
		52 => "011000000110010011100",
		53 => "011000000110010011100",
		54 => "011010100100001110110",
		55 => "011010100100001110110",
		56 => "011010100100001110110",
		57 => "011010100100001010100",
		58 => "011010100100001010100",
		59 => "011010100100001010100",
		60 => "001000111100001010100",
		61 => "001000111100001010100",
		62 => "001000111100001010100",
		63 => "011000001111100010111",
		64 => "011000001111100010111",
		65 => "011000001111100010111",
		66 => "011000101100101010011",
		67 => "011000101100101010011",
		68 => "011000101100101010011",
		69 => "011001100100001110000",
		70 => "011001100100001110000",
		71 => "011001100100001110000",
		72 => "001001011100111010000",
		73 => "001001011100111010000",
		74 => "001001011100111010000",
		75 => "001000011100001010011",
		76 => "001000011100001010011",
		77 => "001000011100001010011",
		78 => "011000000100111010001",
		79 => "011000000100111010001",
		80 => "011000000100111010001",
		81 => "011011011100111010000",
		82 => "011011011100111010000",
		83 => "011011011100111010000",
		84 => "001000100101011010000",
		85 => "001000100101011010000",
		86 => "001000100101011010000",
		87 => "001001011101101010000",
		88 => "001001011101101010000",
		89 => "001001011101101010000",
		90 => "011001000100001110011",
		91 => "011001000100001110011",
		92 => "011001000100001110011",
		93 => "011000000110011011000",
		94 => "011000000110011011000",
		95 => "011000000110011011000",
		96 => "001000011110101010100",
		97 => "001000011110101010100",
		98 => "001000011110101010100",
		99 => "001000010100101011000",
		100 => "001000010100101011000",
		101 => "001000010100101011000",
		102 => "011000001101010010011",
		103 => "011000001101010010011",
		104 => "011000001101010010011",
		105 => "001001111100001010110",
		106 => "001001111100001010110",
		107 => "001001111100001010110",
		108 => "011000000100111110000",
		109 => "011000000100111110000",
		110 => "011000000100111110000",
		111 => "011001100100001110001",
		112 => "011001100100001110001",
		113 => "011001100100001110001",
		114 => "011001100100001110001",
		115 => "011001100100001110001",
		116 => "011001100100001110001",
		117 => "011000000101111010011",
		118 => "011000000101111010011",
		119 => "011000000101111010011",
		120 => "011000001100110110110",
		121 => "011000001100110110110",
		122 => "011000001100110110110",
		123 => "011010100100001010111",
		124 => "011010100100001010111",
		125 => "011010100100001010111",
		126 => "011000001101010010011",
		127 => "011000001101010010011",
		128 => "011000001101010010011",
		129 => "011011000100001010011",
		130 => "011011000100001010011",
		131 => "011011000100001010011",
		132 => "001000011100001010011",
		133 => "001000011100001010011",
		134 => "001000011100001010011",
		135 => "001000111100111010000",
		136 => "001000111100111010000",
		137 => "001000111100111010000",
		138 => "001000111100111010000",
		139 => "001000111100111010000",
		140 => "001000111100111010000",
		141 => "011011100100001110011",
		142 => "011011100100001110011",
		143 => "011011100100001110011",
		144 => "001000011110101010100",
		145 => "001000011110101010100",
		146 => "001000011110101010100",
		147 => "001000010100101011000",
		148 => "001000010100101011000",
		149 => "001000010100101011000",
		150 => "011000001101010010011",
		151 => "011000001101010010011",
		152 => "011000001101010010011",
		153 => "001001111100001010110",
		154 => "001001111100001010110",
		155 => "001001111100001010110",
		156 => "011000000100111110000",
		157 => "011000000100111110000",
		158 => "011000000100111110000",
		159 => "011001100100001110001",
		160 => "011001100100001110001",
		161 => "011001100100001110001",
		162 => "011001100100001110001",
		163 => "011001100100001110001",
		164 => "011001100100001110001",
		165 => "011000000101111010011",
		166 => "011000000101111010011",
		167 => "011000000101111010011",
		168 => "011000001100110110110",
		169 => "011000001100110110110",
		170 => "011000001100110110110",
		171 => "011010100100001010111",
		172 => "011010100100001010111",
		173 => "011010100100001010111",
		174 => "011000001101010010011",
		175 => "011000001101010010011",
		176 => "011000001101010010011",
		177 => "011011000100001010011",
		178 => "011011000100001010011",
		179 => "011011000100001010011",
		180 => "001000011100001010011",
		181 => "001000011100001010011",
		182 => "001000011100001010011",
		183 => "001000111100111010000",
		184 => "001000111100111010000",
		185 => "001000111100111010000",
		186 => "001000111100111010000",
		187 => "001000111100111010000",
		188 => "001000111100111010000",
		189 => "011011100100001110011",
		190 => "011011100100001110011",
		191 => "011011100100001110011",
		192 => "011100000100001010011",
		193 => "011100000100001010011",
		194 => "011100000100001010011",
		195 => "011000000101111011000",
		196 => "011000000101111011000",
		197 => "011000000101111011000",
		198 => "001011011100001110010",
		199 => "001011011100001110010",
		200 => "001011011100001110010",
		201 => "011000000101101010011",
		202 => "011000000101101010011",
		203 => "011000000101101010011",
		204 => "011100000100001111001",
		205 => "011100000100001111001",
		206 => "011100000100001111001",
		207 => "001000111100001010011",
		208 => "001000111100001010011",
		209 => "001000111100001010011",
		210 => "001000000100101010110",
		211 => "001000000100101010110",
		212 => "001000000100101010110",
		213 => "001001100101101010000",
		214 => "001001100101101010000",
		215 => "001001100101101010000",
		216 => "011100000100001010011",
		217 => "011100000100001010011",
		218 => "011100000100001010011",
		219 => "011000000101111011000",
		220 => "011000000101111011000",
		221 => "011000000101111011000",
		222 => "001011011100001110010",
		223 => "001011011100001110010",
		224 => "001011011100001110010",
		225 => "011000000101101010011",
		226 => "011000000101101010011",
		227 => "011000000101101010011",
		228 => "011100000100001111001",
		229 => "011100000100001111001",
		230 => "011100000100001111001",
		231 => "001000111100001010011",
		232 => "001000111100001010011",
		233 => "001000111100001010011",
		234 => "001000000100101010110",
		235 => "001000000100101010110",
		236 => "001000000100101010110",
		237 => "001001100101101010000",
		238 => "001001100101101010000",
		239 => "001001100101101010000",
		240 => "011100000100001010011",
		241 => "011100000100001010011",
		242 => "011100000100001010011",
		243 => "011000000101111011000",
		244 => "011000000101111011000",
		245 => "011000000101111011000",
		246 => "001011011100001110010",
		247 => "001011011100001110010",
		248 => "001011011100001110010",
		249 => "011000000101101010011",
		250 => "011000000101101010011",
		251 => "011000000101101010011",
		252 => "011100000100001111001",
		253 => "011100000100001111001",
		254 => "011100000100001111001",
		255 => "001000111100001010011",
		256 => "001000111100001010011",
		257 => "001000111100001010011",
		258 => "001000000100101010110",
		259 => "001000000100101010110",
		260 => "001000000100101010110",
		261 => "001001100101101010000",
		262 => "001001100101101010000",
		263 => "001001100101101010000",
		264 => "011100000100001010011",
		265 => "011100000100001010011",
		266 => "011100000100001010011",
		267 => "011000000101111011000",
		268 => "011000000101111011000",
		269 => "011000000101111011000",
		270 => "001011011100001110010",
		271 => "001011011100001110010",
		272 => "001011011100001110010",
		273 => "011000000101101010011",
		274 => "011000000101101010011",
		275 => "011000000101101010011",
		276 => "011100000100001111001",
		277 => "011100000100001111001",
		278 => "011100000100001111001",
		279 => "001000111100001010011",
		280 => "001000111100001010011",
		281 => "001000111100001010011",
		282 => "001000000100101010110",
		283 => "001000000100101010110",
		284 => "001000000100101010110",
		285 => "001001100101101010000",
		286 => "001001100101101010000",
		287 => "001001100101101010000",
		288 => "011000001110100010101",
		289 => "011000001110100010101",
		290 => "011000001110100010101",
		291 => "011000111100001010011",
		292 => "011000111100001010011",
		293 => "011000111100001010011",
		294 => "011000001110100010101",
		295 => "011000001110100010101",
		296 => "011000001110100010101",
		297 => "011001100100001110001",
		298 => "011001100100001110001",
		299 => "011001100100001110001",
		300 => "011000001110100010101",
		301 => "011000001110100010101",
		302 => "011000001110100010101",
		303 => "011000111100001010011",
		304 => "011000111100001010011",
		305 => "011000111100001010011",
		306 => "011000001110100010101",
		307 => "011000001110100010101",
		308 => "011000001110100010101",
		309 => "011001100100001110001",
		310 => "011001100100001110001",
		311 => "011001100100001110001",
		312 => "011000001110100010101",
		313 => "011000001110100010101",
		314 => "011000001110100010101",
		315 => "011000111100001010011",
		316 => "011000111100001010011",
		317 => "011000111100001010011",
		318 => "011000001110100010101",
		319 => "011000001110100010101",
		320 => "011000001110100010101",
		321 => "011001100100001110001",
		322 => "011001100100001110001",
		323 => "011001100100001110001",
		324 => "011000001110100010101",
		325 => "011000001110100010101",
		326 => "011000001110100010101",
		327 => "011000111100001010011",
		328 => "011000111100001010011",
		329 => "011000111100001010011",
		330 => "011000001110100010101",
		331 => "011000001110100010101",
		332 => "011000001110100010101",
		333 => "011001100100001110001",
		334 => "011001100100001110001",
		335 => "011001100100001110001",
		336 => "011000001110100010101",
		337 => "011000001110100010101",
		338 => "011000001110100010101",
		339 => "011000111100001010011",
		340 => "011000111100001010011",
		341 => "011000111100001010011",
		342 => "011000001110100010101",
		343 => "011000001110100010101",
		344 => "011000001110100010101",
		345 => "011001100100001110001",
		346 => "011001100100001110001",
		347 => "011001100100001110001",
		348 => "011000001110100010101",
		349 => "011000001110100010101",
		350 => "011000001110100010101",
		351 => "011000111100001010011",
		352 => "011000111100001010011",
		353 => "011000111100001010011",
		354 => "011000001110100010101",
		355 => "011000001110100010101",
		356 => "011000001110100010101",
		357 => "011001100100001110001",
		358 => "011001100100001110001",
		359 => "011001100100001110001",
		360 => "011000001110100010101",
		361 => "011000001110100010101",
		362 => "011000001110100010101",
		363 => "011000111100001010011",
		364 => "011000111100001010011",
		365 => "011000111100001010011",
		366 => "011000001110100010101",
		367 => "011000001110100010101",
		368 => "011000001110100010101",
		369 => "011001100100001110001",
		370 => "011001100100001110001",
		371 => "011001100100001110001",
		372 => "011000001110100010101",
		373 => "011000001110100010101",
		374 => "011000001110100010101",
		375 => "011000111100001010011",
		376 => "011000111100001010011",
		377 => "011000111100001010011",
		378 => "011000001110100010101",
		379 => "011000001110100010101",
		380 => "011000001110100010101",
		381 => "011001100100001110001",
		382 => "011001100100001110001",
		383 => "011001100100001110001",
		384 => "011001011101001010000",
		385 => "011001011101001010000",
		386 => "011001011101001010000",
		387 => "011010000100001010010",
		388 => "011010000100001010010",
		389 => "011010000100001010010",
		390 => "011001011101001010000",
		391 => "011001011101001010000",
		392 => "011001011101001010000",
		393 => "011010000100001010010",
		394 => "011010000100001010010",
		395 => "011010000100001010010",
		396 => "011001011101001010000",
		397 => "011001011101001010000",
		398 => "011001011101001010000",
		399 => "011010000100001010010",
		400 => "011010000100001010010",
		401 => "011010000100001010010",
		402 => "011001011101001010000",
		403 => "011001011101001010000",
		404 => "011001011101001010000",
		405 => "011010000100001010010",
		406 => "011010000100001010010",
		407 => "011010000100001010010",
		408 => "011001011101001010000",
		409 => "011001011101001010000",
		410 => "011001011101001010000",
		411 => "011010000100001010010",
		412 => "011010000100001010010",
		413 => "011010000100001010010",
		414 => "011001011101001010000",
		415 => "011001011101001010000",
		416 => "011001011101001010000",
		417 => "011010000100001010010",
		418 => "011010000100001010010",
		419 => "011010000100001010010",
		420 => "011001011101001010000",
		421 => "011001011101001010000",
		422 => "011001011101001010000",
		423 => "011010000100001010010",
		424 => "011010000100001010010",
		425 => "011010000100001010010",
		426 => "011001011101001010000",
		427 => "011001011101001010000",
		428 => "011001011101001010000",
		429 => "011010000100001010010",
		430 => "011010000100001010010",
		431 => "011010000100001010010",
		432 => "011001011101001010000",
		433 => "011001011101001010000",
		434 => "011001011101001010000",
		435 => "011010000100001010010",
		436 => "011010000100001010010",
		437 => "011010000100001010010",
		438 => "011001011101001010000",
		439 => "011001011101001010000",
		440 => "011001011101001010000",
		441 => "011010000100001010010",
		442 => "011010000100001010010",
		443 => "011010000100001010010",
		444 => "011001011101001010000",
		445 => "011001011101001010000",
		446 => "011001011101001010000",
		447 => "011010000100001010010",
		448 => "011010000100001010010",
		449 => "011010000100001010010",
		450 => "011001011101001010000",
		451 => "011001011101001010000",
		452 => "011001011101001010000",
		453 => "011010000100001010010",
		454 => "011010000100001010010",
		455 => "011010000100001010010",
		456 => "011001011101001010000",
		457 => "011001011101001010000",
		458 => "011001011101001010000",
		459 => "011010000100001010010",
		460 => "011010000100001010010",
		461 => "011010000100001010010",
		462 => "011001011101001010000",
		463 => "011001011101001010000",
		464 => "011001011101001010000",
		465 => "011010000100001010010",
		466 => "011010000100001010010",
		467 => "011010000100001010010",
		468 => "011001011101001010000",
		469 => "011001011101001010000",
		470 => "011001011101001010000",
		471 => "011010000100001010010",
		472 => "011010000100001010010",
		473 => "011010000100001010010",
		474 => "011001011101001010000",
		475 => "011001011101001010000",
		476 => "011001011101001010000",
		477 => "011010000100001010010",
		478 => "011010000100001010010",
		479 => "011010000100001010010",
		480 => "111011010100001010011",
		481 => "111011010100001010011",
		482 => "111011010100001010011",
		483 => "111011010100001010011",
		484 => "111011010100001010011",
		485 => "111011010100001010011",
		486 => "111011010100001010011",
		487 => "111011010100001010011",
		488 => "111011010100001010011",
		489 => "111011010100001010011",
		490 => "111011010100001010011",
		491 => "111011010100001010011",
		492 => "111011010100001010011",
		493 => "111011010100001010011",
		494 => "111011010100001010011",
		495 => "111011010100001010011",
		496 => "111011010100001010011",
		497 => "111011010100001010011",
		498 => "111011010100001010011",
		499 => "111011010100001010011",
		500 => "111011010100001010011",
		501 => "111011010100001010011",
		502 => "111011010100001010011",
		503 => "111011010100001010011",
		504 => "111011010100001010011",
		505 => "111011010100001010011",
		506 => "111011010100001010011",
		507 => "111011010100001010011",
		508 => "111011010100001010011",
		509 => "111011010100001010011",
		510 => "111011010100001010011",
		511 => "111011010100001010011",
		512 => "111011010100001010011",
		513 => "111011010100001010011",
		514 => "111011010100001010011",
		515 => "111011010100001010011",
		516 => "111011010100001010011",
		517 => "111011010100001010011",
		518 => "111011010100001010011",
		519 => "111011010100001010011",
		520 => "111011010100001010011",
		521 => "111011010100001010011",
		522 => "111011010100001010011",
		523 => "111011010100001010011",
		524 => "111011010100001010011",
		525 => "111011010100001010011",
		526 => "111011010100001010011",
		527 => "111011010100001010011",
		528 => "111011010100001010011",
		529 => "111011010100001010011",
		530 => "111011010100001010011",
		531 => "111011010100001010011",
		532 => "111011010100001010011",
		533 => "111011010100001010011",
		534 => "111011010100001010011",
		535 => "111011010100001010011",
		536 => "111011010100001010011",
		537 => "111011010100001010011",
		538 => "111011010100001010011",
		539 => "111011010100001010011",
		540 => "111011010100001010011",
		541 => "111011010100001010011",
		542 => "111011010100001010011",
		543 => "111011010100001010011",
		544 => "111011010100001010011",
		545 => "111011010100001010011",
		546 => "111011010100001010011",
		547 => "111011010100001010011",
		548 => "111011010100001010011",
		549 => "111011010100001010011",
		550 => "111011010100001010011",
		551 => "111011010100001010011",
		552 => "111011010100001010011",
		553 => "111011010100001010011",
		554 => "111011010100001010011",
		555 => "111011010100001010011",
		556 => "111011010100001010011",
		557 => "111011010100001010011",
		558 => "111011010100001010011",
		559 => "111011010100001010011",
		560 => "111011010100001010011",
		561 => "111011010100001010011",
		562 => "111011010100001010011",
		563 => "111011010100001010011",
		564 => "111011010100001010011",
		565 => "111011010100001010011",
		566 => "111011010100001010011",
		567 => "111011010100001010011",
		568 => "111011010100001010011",
		569 => "111011010100001010011",
		570 => "111011010100001010011",
		571 => "111011010100001010011",
		572 => "111011010100001010011",
		573 => "111011010100001010011",
		574 => "111011010100001010011",
		575 => "111011010100001010011",
		576 => "011011000100001110011",
		577 => "011011000100001110011",
		578 => "011011000100001110011",
		579 => "011011000100001110011",
		580 => "011011000100001110011",
		581 => "011011000100001110011",
		582 => "011011000100001110011",
		583 => "011011000100001110011",
		584 => "011011000100001110011",
		585 => "011011000100001110011",
		586 => "011011000100001110011",
		587 => "011011000100001110011",
		588 => "011011000100001110011",
		589 => "011011000100001110011",
		590 => "011011000100001110011",
		591 => "011011000100001110011",
		592 => "011011000100001110011",
		593 => "011011000100001110011",
		594 => "011011000100001110011",
		595 => "011011000100001110011",
		596 => "011011000100001110011",
		597 => "011011000100001110011",
		598 => "011011000100001110011",
		599 => "011011000100001110011",
		600 => "011011000100001110011",
		601 => "011011000100001110011",
		602 => "011011000100001110011",
		603 => "011011000100001110011",
		604 => "011011000100001110011",
		605 => "011011000100001110011",
		606 => "011011000100001110011",
		607 => "011011000100001110011",
		608 => "011011000100001110011",
		609 => "011011000100001110011",
		610 => "011011000100001110011",
		611 => "011011000100001110011",
		612 => "011011000100001110011",
		613 => "011011000100001110011",
		614 => "011011000100001110011",
		615 => "011011000100001110011",
		616 => "011011000100001110011",
		617 => "011011000100001110011",
		618 => "011011000100001110011",
		619 => "011011000100001110011",
		620 => "011011000100001110011",
		621 => "011011000100001110011",
		622 => "011011000100001110011",
		623 => "011011000100001110011",
		624 => "011011000100001110011",
		625 => "011011000100001110011",
		626 => "011011000100001110011",
		627 => "011011000100001110011",
		628 => "011011000100001110011",
		629 => "011011000100001110011",
		630 => "011011000100001110011",
		631 => "011011000100001110011",
		632 => "011011000100001110011",
		633 => "011011000100001110011",
		634 => "011011000100001110011",
		635 => "011011000100001110011",
		636 => "011011000100001110011",
		637 => "011011000100001110011",
		638 => "011011000100001110011",
		639 => "011011000100001110011",
		640 => "011011000100001110011",
		641 => "011011000100001110011",
		642 => "011011000100001110011",
		643 => "011011000100001110011",
		644 => "011011000100001110011",
		645 => "011011000100001110011",
		646 => "011011000100001110011",
		647 => "011011000100001110011",
		648 => "011011000100001110011",
		649 => "011011000100001110011",
		650 => "011011000100001110011",
		651 => "011011000100001110011",
		652 => "011011000100001110011",
		653 => "011011000100001110011",
		654 => "011011000100001110011",
		655 => "011011000100001110011",
		656 => "011011000100001110011",
		657 => "011011000100001110011",
		658 => "011011000100001110011",
		659 => "011011000100001110011",
		660 => "011011000100001110011",
		661 => "011011000100001110011",
		662 => "011011000100001110011",
		663 => "011011000100001110011",
		664 => "011011000100001110011",
		665 => "011011000100001110011",
		666 => "011011000100001110011",
		667 => "011011000100001110011",
		668 => "011011000100001110011",
		669 => "011011000100001110011",
		670 => "011011000100001110011",
		671 => "011011000100001110011",
		672 => "011000101100100010101",
		673 => "011000101100100010101",
		674 => "011000101100100010101",
		675 => "011000101100100010101",
		676 => "011000101100100010101",
		677 => "011000101100100010101",
		678 => "011000101100100010101",
		679 => "011000101100100010101",
		680 => "011000101100100010101",
		681 => "011000101100100010101",
		682 => "011000101100100010101",
		683 => "011000101100100010101",
		684 => "011000101100100010101",
		685 => "011000101100100010101",
		686 => "011000101100100010101",
		687 => "011000101100100010101",
		688 => "011000101100100010101",
		689 => "011000101100100010101",
		690 => "011000101100100010101",
		691 => "011000101100100010101",
		692 => "011000101100100010101",
		693 => "011000101100100010101",
		694 => "011000101100100010101",
		695 => "011000101100100010101",
		696 => "011000101100100010101",
		697 => "011000101100100010101",
		698 => "011000101100100010101",
		699 => "011000101100100010101",
		700 => "011000101100100010101",
		701 => "011000101100100010101",
		702 => "011000101100100010101",
		703 => "011000101100100010101",
		704 => "011000101100100010101",
		705 => "011000101100100010101",
		706 => "011000101100100010101",
		707 => "011000101100100010101",
		708 => "011000101100100010101",
		709 => "011000101100100010101",
		710 => "011000101100100010101",
		711 => "011000101100100010101",
		712 => "011000101100100010101",
		713 => "011000101100100010101",
		714 => "011000101100100010101",
		715 => "011000101100100010101",
		716 => "011000101100100010101",
		717 => "011000101100100010101",
		718 => "011000101100100010101",
		719 => "011000101100100010101",
		720 => "011000101100100010101",
		721 => "011000101100100010101",
		722 => "011000101100100010101",
		723 => "011000101100100010101",
		724 => "011000101100100010101",
		725 => "011000101100100010101",
		726 => "011000101100100010101",
		727 => "011000101100100010101",
		728 => "011000101100100010101",
		729 => "011000101100100010101",
		730 => "011000101100100010101",
		731 => "011000101100100010101",
		732 => "011000101100100010101",
		733 => "011000101100100010101",
		734 => "011000101100100010101",
		735 => "011000101100100010101",
		736 => "011000101100100010101",
		737 => "011000101100100010101",
		738 => "011000101100100010101",
		739 => "011000101100100010101",
		740 => "011000101100100010101",
		741 => "011000101100100010101",
		742 => "011000101100100010101",
		743 => "011000101100100010101",
		744 => "011000101100100010101",
		745 => "011000101100100010101",
		746 => "011000101100100010101",
		747 => "011000101100100010101",
		748 => "011000101100100010101",
		749 => "011000101100100010101",
		750 => "011000101100100010101",
		751 => "011000101100100010101",
		752 => "011000101100100010101",
		753 => "011000101100100010101",
		754 => "011000101100100010101",
		755 => "011000101100100010101",
		756 => "011000101100100010101",
		757 => "011000101100100010101",
		758 => "011000101100100010101",
		759 => "011000101100100010101",
		760 => "011000101100100010101",
		761 => "011000101100100010101",
		762 => "011000101100100010101",
		763 => "011000101100100010101",
		764 => "011000101100100010101",
		765 => "011000101100100010101",
		766 => "011000101100100010101",
		767 => "011000101100100010101",
		768 => "011000101100100110010",
		769 => "011000101100100110010",
		770 => "011000101100100110010",
		771 => "011000101100100110010",
		772 => "011000101100100110010",
		773 => "011000101100100110010",
		774 => "011000101100100110010",
		775 => "011000101100100110010",
		776 => "011000101100100110010",
		777 => "011000101100100110010",
		778 => "011000101100100110010",
		779 => "011000101100100110010",
		780 => "011000101100100110010",
		781 => "011000101100100110010",
		782 => "011000101100100110010",
		783 => "011000101100100110010",
		784 => "011000101100100110010",
		785 => "011000101100100110010",
		786 => "011000101100100110010",
		787 => "011000101100100110010",
		788 => "011000101100100110010",
		789 => "011000101100100110010",
		790 => "011000101100100110010",
		791 => "011000101100100110010",
		792 => "011000101100100110010",
		793 => "011000101100100110010",
		794 => "011000101100100110010",
		795 => "011000101100100110010",
		796 => "011000101100100110010",
		797 => "011000101100100110010",
		798 => "011000101100100110010",
		799 => "011000101100100110010",
		800 => "011000101100100110010",
		801 => "011000101100100110010",
		802 => "011000101100100110010",
		803 => "011000101100100110010",
		804 => "011000101100100110010",
		805 => "011000101100100110010",
		806 => "011000101100100110010",
		807 => "011000101100100110010",
		808 => "011000101100100110010",
		809 => "011000101100100110010",
		810 => "011000101100100110010",
		811 => "011000101100100110010",
		812 => "011000101100100110010",
		813 => "011000101100100110010",
		814 => "011000101100100110010",
		815 => "011000101100100110010",
		816 => "011000101100100110010",
		817 => "011000101100100110010",
		818 => "011000101100100110010",
		819 => "011000101100100110010",
		820 => "011000101100100110010",
		821 => "011000101100100110010",
		822 => "011000101100100110010",
		823 => "011000101100100110010",
		824 => "011000101100100110010",
		825 => "011000101100100110010",
		826 => "011000101100100110010",
		827 => "011000101100100110010",
		828 => "011000101100100110010",
		829 => "011000101100100110010",
		830 => "011000101100100110010",
		831 => "011000101100100110010",
		832 => "011000101100100110010",
		833 => "011000101100100110010",
		834 => "011000101100100110010",
		835 => "011000101100100110010",
		836 => "011000101100100110010",
		837 => "011000101100100110010",
		838 => "011000101100100110010",
		839 => "011000101100100110010",
		840 => "011000101100100110010",
		841 => "011000101100100110010",
		842 => "011000101100100110010",
		843 => "011000101100100110010",
		844 => "011000101100100110010",
		845 => "011000101100100110010",
		846 => "011000101100100110010",
		847 => "011000101100100110010",
		848 => "011000101100100110010",
		849 => "011000101100100110010",
		850 => "011000101100100110010",
		851 => "011000101100100110010",
		852 => "011000101100100110010",
		853 => "011000101100100110010",
		854 => "011000101100100110010",
		855 => "011000101100100110010",
		856 => "011000101100100110010",
		857 => "011000101100100110010",
		858 => "011000101100100110010",
		859 => "011000101100100110010",
		860 => "011000101100100110010",
		861 => "011000101100100110010",
		862 => "011000101100100110010",
		863 => "011000101100100110010");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;