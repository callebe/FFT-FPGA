library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT1024p_5 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT1024p_5;

architecture Behavioral of ROMFFT1024p_5 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 6 
	constant ROM_tb : ROM := (
		0 => "001101111110111010000",
		1 => "001101111110111010000",
		2 => "001101111110111010000",
		3 => "001011011100001011001",
		4 => "001011011100001011001",
		5 => "001011011100001011001",
		6 => "001010000110001110000",
		7 => "001010000110001110000",
		8 => "001010000110001110000",
		9 => "011011100100001010011",
		10 => "011011100100001010011",
		11 => "011011100100001010011",
		12 => "011011011100001010101",
		13 => "011011011100001010101",
		14 => "011011011100001010101",
		15 => "011000001110100010101",
		16 => "011000001110100010101",
		17 => "011000001110100010101",
		18 => "001010011100001010101",
		19 => "001010011100001010101",
		20 => "001010011100001010101",
		21 => "001001011100001010111",
		22 => "001001011100001010111",
		23 => "001001011100001010111",
		24 => "011010000100001010001",
		25 => "011010000100001010001",
		26 => "011010000100001010001",
		27 => "011001011101001010000",
		28 => "011001011101001010000",
		29 => "011001011101001010000",
		30 => "011000000100111110001",
		31 => "011000000100111110001",
		32 => "011000000100111110001",
		33 => "001000111100011110010",
		34 => "001000111100011110010",
		35 => "001000111100011110010",
		36 => "011000101100101010011",
		37 => "011000101100101010011",
		38 => "011000101100101010011",
		39 => "011000110100011010011",
		40 => "011000110100011010011",
		41 => "011000110100011010011",
		42 => "011000000100111010000",
		43 => "011000000100111010000",
		44 => "011000000100111010000",
		45 => "011000011100111010000",
		46 => "011000011100111010000",
		47 => "011000011100111010000",
		48 => "001001011100111010000",
		49 => "001001011100111010000",
		50 => "001001011100111010000",
		51 => "001000100100111110001",
		52 => "001000100100111110001",
		53 => "001000100100111110001",
		54 => "011000011100111010000",
		55 => "011000011100111010000",
		56 => "011000011100111010000",
		57 => "011001001100111110000",
		58 => "011001001100111110000",
		59 => "011001001100111110000",
		60 => "011000000100111010001",
		61 => "011000000100111010001",
		62 => "011000000100111010001",
		63 => "011001011100001010100",
		64 => "011001011100001010100",
		65 => "011001011100001010100",
		66 => "001011011100001010011",
		67 => "001011011100001010011",
		68 => "001011011100001010011",
		69 => "011000000100111010001",
		70 => "011000000100111010001",
		71 => "011000000100111010001",
		72 => "001000011100011110101",
		73 => "001000011100011110101",
		74 => "001000011100011110101",
		75 => "011010011100001010101",
		76 => "011010011100001010101",
		77 => "011010011100001010101",
		78 => "011000000101101010010",
		79 => "011000000101101010010",
		80 => "011000000101101010010",
		81 => "001000000100111110010",
		82 => "001000000100111110010",
		83 => "001000000100111110010",
		84 => "011000101100101010011",
		85 => "011000101100101010011",
		86 => "011000101100101010011",
		87 => "011000001111010010111",
		88 => "011000001111010010111",
		89 => "011000001111010010111",
		90 => "011000000110011011000",
		91 => "011000000110011011000",
		92 => "011000000110011011000",
		93 => "011000011110101011000",
		94 => "011000011110101011000",
		95 => "011000011110101011000",
		96 => "001000011110101010100",
		97 => "001000011110101010100",
		98 => "001000011110101010100",
		99 => "011001111101111010000",
		100 => "011001111101111010000",
		101 => "011001111101111010000",
		102 => "001000010100101011000",
		103 => "001000010100101011000",
		104 => "001000010100101011000",
		105 => "011001001100111010000",
		106 => "011001001100111010000",
		107 => "011001001100111010000",
		108 => "011000001101010010011",
		109 => "011000001101010010011",
		110 => "011000001101010010011",
		111 => "011000111101001010000",
		112 => "011000111101001010000",
		113 => "011000111101001010000",
		114 => "001001111100001010110",
		115 => "001001111100001010110",
		116 => "001001111100001010110",
		117 => "001001011100001010011",
		118 => "001001011100001010011",
		119 => "001001011100001010011",
		120 => "011000000100111110000",
		121 => "011000000100111110000",
		122 => "011000000100111110000",
		123 => "001010011100011110010",
		124 => "001010011100011110010",
		125 => "001010011100011110010",
		126 => "011001100100001110001",
		127 => "011001100100001110001",
		128 => "011001100100001110001",
		129 => "011000000101001010100",
		130 => "011000000101001010100",
		131 => "011000000101001010100",
		132 => "011001100100001110001",
		133 => "011001100100001110001",
		134 => "011001100100001110001",
		135 => "011000000101101010010",
		136 => "011000000101101010010",
		137 => "011000000101101010010",
		138 => "011000000101111010011",
		139 => "011000000101111010011",
		140 => "011000000101111010011",
		141 => "011100001110011110000",
		142 => "011100001110011110000",
		143 => "011100001110011110000",
		144 => "011000001100110110110",
		145 => "011000001100110110110",
		146 => "011000001100110110110",
		147 => "011011100100001010011",
		148 => "011011100100001010011",
		149 => "011011100100001010011",
		150 => "011010100100001010111",
		151 => "011010100100001010111",
		152 => "011010100100001010111",
		153 => "011001100100011110000",
		154 => "011001100100011110000",
		155 => "011001100100011110000",
		156 => "011000001101010010011",
		157 => "011000001101010010011",
		158 => "011000001101010010011",
		159 => "011000111101001010000",
		160 => "011000111101001010000",
		161 => "011000111101001010000",
		162 => "011011000100001010011",
		163 => "011011000100001010011",
		164 => "011011000100001010011",
		165 => "011001100100001010010",
		166 => "011001100100001010010",
		167 => "011001100100001010010",
		168 => "001000011100001010011",
		169 => "001000011100001010011",
		170 => "001000011100001010011",
		171 => "011001000100001010100",
		172 => "011001000100001010100",
		173 => "011001000100001010100",
		174 => "001000111100111010000",
		175 => "001000111100111010000",
		176 => "001000111100111010000",
		177 => "011010000100001110100",
		178 => "011010000100001110100",
		179 => "011010000100001110100",
		180 => "001000111100111010000",
		181 => "001000111100111010000",
		182 => "001000111100111010000",
		183 => "011000000101101010010",
		184 => "011000000101101010010",
		185 => "011000000101101010010",
		186 => "011011100100001110011",
		187 => "011011100100001110011",
		188 => "011011100100001110011",
		189 => "001000011110001111001",
		190 => "001000011110001111001",
		191 => "001000011110001111001",
		192 => "011100000100001010011",
		193 => "011100000100001010011",
		194 => "011100000100001010011",
		195 => "001001011100001010101",
		196 => "001001011100001010101",
		197 => "001001011100001010101",
		198 => "011000000101111011000",
		199 => "011000000101111011000",
		200 => "011000000101111011000",
		201 => "001010011100011110010",
		202 => "001010011100011110010",
		203 => "001010011100011110010",
		204 => "001011011100001110010",
		205 => "001011011100001110010",
		206 => "001011011100001110010",
		207 => "011000001101100010011",
		208 => "011000001101100010011",
		209 => "011000001101100010011",
		210 => "011000000101101010011",
		211 => "011000000101101010011",
		212 => "011000000101101010011",
		213 => "011000011110001010110",
		214 => "011000011110001010110",
		215 => "011000011110001010110",
		216 => "011100000100001111001",
		217 => "011100000100001111001",
		218 => "011100000100001111001",
		219 => "011010100100001010010",
		220 => "011010100100001010010",
		221 => "011010100100001010010",
		222 => "001000111100001010011",
		223 => "001000111100001010011",
		224 => "001000111100001010011",
		225 => "011001000100001010100",
		226 => "011001000100001010100",
		227 => "011001000100001010100",
		228 => "001000000100101010110",
		229 => "001000000100101010110",
		230 => "001000000100101010110",
		231 => "011000001101100010011",
		232 => "011000001101100010011",
		233 => "011000001101100010011",
		234 => "001001100101101010000",
		235 => "001001100101101010000",
		236 => "001001100101101010000",
		237 => "011100000101101010000",
		238 => "011100000101101010000",
		239 => "011100000101101010000",
		240 => "011100000100001010011",
		241 => "011100000100001010011",
		242 => "011100000100001010011",
		243 => "001001011100001010101",
		244 => "001001011100001010101",
		245 => "001001011100001010101",
		246 => "011000000101111011000",
		247 => "011000000101111011000",
		248 => "011000000101111011000",
		249 => "001010011100011110010",
		250 => "001010011100011110010",
		251 => "001010011100011110010",
		252 => "001011011100001110010",
		253 => "001011011100001110010",
		254 => "001011011100001110010",
		255 => "011000001101100010011",
		256 => "011000001101100010011",
		257 => "011000001101100010011",
		258 => "011000000101101010011",
		259 => "011000000101101010011",
		260 => "011000000101101010011",
		261 => "011000011110001010110",
		262 => "011000011110001010110",
		263 => "011000011110001010110",
		264 => "011100000100001111001",
		265 => "011100000100001111001",
		266 => "011100000100001111001",
		267 => "011010100100001010010",
		268 => "011010100100001010010",
		269 => "011010100100001010010",
		270 => "001000111100001010011",
		271 => "001000111100001010011",
		272 => "001000111100001010011",
		273 => "011001000100001010100",
		274 => "011001000100001010100",
		275 => "011001000100001010100",
		276 => "001000000100101010110",
		277 => "001000000100101010110",
		278 => "001000000100101010110",
		279 => "011000001101100010011",
		280 => "011000001101100010011",
		281 => "011000001101100010011",
		282 => "001001100101101010000",
		283 => "001001100101101010000",
		284 => "001001100101101010000",
		285 => "011100000101101010000",
		286 => "011100000101101010000",
		287 => "011100000101101010000",
		288 => "011000001110100010101",
		289 => "011000001110100010101",
		290 => "011000001110100010101",
		291 => "001001111100001010110",
		292 => "001001111100001010110",
		293 => "001001111100001010110",
		294 => "011000111100001010011",
		295 => "011000111100001010011",
		296 => "011000111100001010011",
		297 => "011000010100111010110",
		298 => "011000010100111010110",
		299 => "011000010100111010110",
		300 => "011000001110100010101",
		301 => "011000001110100010101",
		302 => "011000001110100010101",
		303 => "011011000100001010011",
		304 => "011011000100001010011",
		305 => "011011000100001010011",
		306 => "011001100100001110001",
		307 => "011001100100001110001",
		308 => "011001100100001110001",
		309 => "011000000101110011001",
		310 => "011000000101110011001",
		311 => "011000000101110011001",
		312 => "011000001110100010101",
		313 => "011000001110100010101",
		314 => "011000001110100010101",
		315 => "001001111100001010110",
		316 => "001001111100001010110",
		317 => "001001111100001010110",
		318 => "011000111100001010011",
		319 => "011000111100001010011",
		320 => "011000111100001010011",
		321 => "011000010100111010110",
		322 => "011000010100111010110",
		323 => "011000010100111010110",
		324 => "011000001110100010101",
		325 => "011000001110100010101",
		326 => "011000001110100010101",
		327 => "011011000100001010011",
		328 => "011011000100001010011",
		329 => "011011000100001010011",
		330 => "011001100100001110001",
		331 => "011001100100001110001",
		332 => "011001100100001110001",
		333 => "011000000101110011001",
		334 => "011000000101110011001",
		335 => "011000000101110011001",
		336 => "011000001110100010101",
		337 => "011000001110100010101",
		338 => "011000001110100010101",
		339 => "001001111100001010110",
		340 => "001001111100001010110",
		341 => "001001111100001010110",
		342 => "011000111100001010011",
		343 => "011000111100001010011",
		344 => "011000111100001010011",
		345 => "011000010100111010110",
		346 => "011000010100111010110",
		347 => "011000010100111010110",
		348 => "011000001110100010101",
		349 => "011000001110100010101",
		350 => "011000001110100010101",
		351 => "011011000100001010011",
		352 => "011011000100001010011",
		353 => "011011000100001010011",
		354 => "011001100100001110001",
		355 => "011001100100001110001",
		356 => "011001100100001110001",
		357 => "011000000101110011001",
		358 => "011000000101110011001",
		359 => "011000000101110011001",
		360 => "011000001110100010101",
		361 => "011000001110100010101",
		362 => "011000001110100010101",
		363 => "001001111100001010110",
		364 => "001001111100001010110",
		365 => "001001111100001010110",
		366 => "011000111100001010011",
		367 => "011000111100001010011",
		368 => "011000111100001010011",
		369 => "011000010100111010110",
		370 => "011000010100111010110",
		371 => "011000010100111010110",
		372 => "011000001110100010101",
		373 => "011000001110100010101",
		374 => "011000001110100010101",
		375 => "011011000100001010011",
		376 => "011011000100001010011",
		377 => "011011000100001010011",
		378 => "011001100100001110001",
		379 => "011001100100001110001",
		380 => "011001100100001110001",
		381 => "011000000101110011001",
		382 => "011000000101110011001",
		383 => "011000000101110011001",
		384 => "011001011101001010000",
		385 => "011001011101001010000",
		386 => "011001011101001010000",
		387 => "011000000101011010101",
		388 => "011000000101011010101",
		389 => "011000000101011010101",
		390 => "011010000100001010010",
		391 => "011010000100001010010",
		392 => "011010000100001010010",
		393 => "011000000101011010101",
		394 => "011000000101011010101",
		395 => "011000000101011010101",
		396 => "011001011101001010000",
		397 => "011001011101001010000",
		398 => "011001011101001010000",
		399 => "011000000101011010101",
		400 => "011000000101011010101",
		401 => "011000000101011010101",
		402 => "011010000100001010010",
		403 => "011010000100001010010",
		404 => "011010000100001010010",
		405 => "011000000101011010101",
		406 => "011000000101011010101",
		407 => "011000000101011010101",
		408 => "011001011101001010000",
		409 => "011001011101001010000",
		410 => "011001011101001010000",
		411 => "011000000101011010101",
		412 => "011000000101011010101",
		413 => "011000000101011010101",
		414 => "011010000100001010010",
		415 => "011010000100001010010",
		416 => "011010000100001010010",
		417 => "011000000101011010101",
		418 => "011000000101011010101",
		419 => "011000000101011010101",
		420 => "011001011101001010000",
		421 => "011001011101001010000",
		422 => "011001011101001010000",
		423 => "011000000101011010101",
		424 => "011000000101011010101",
		425 => "011000000101011010101",
		426 => "011010000100001010010",
		427 => "011010000100001010010",
		428 => "011010000100001010010",
		429 => "011000000101011010101",
		430 => "011000000101011010101",
		431 => "011000000101011010101",
		432 => "011001011101001010000",
		433 => "011001011101001010000",
		434 => "011001011101001010000",
		435 => "011000000101011010101",
		436 => "011000000101011010101",
		437 => "011000000101011010101",
		438 => "011010000100001010010",
		439 => "011010000100001010010",
		440 => "011010000100001010010",
		441 => "011000000101011010101",
		442 => "011000000101011010101",
		443 => "011000000101011010101",
		444 => "011001011101001010000",
		445 => "011001011101001010000",
		446 => "011001011101001010000",
		447 => "011000000101011010101",
		448 => "011000000101011010101",
		449 => "011000000101011010101",
		450 => "011010000100001010010",
		451 => "011010000100001010010",
		452 => "011010000100001010010",
		453 => "011000000101011010101",
		454 => "011000000101011010101",
		455 => "011000000101011010101",
		456 => "011001011101001010000",
		457 => "011001011101001010000",
		458 => "011001011101001010000",
		459 => "011000000101011010101",
		460 => "011000000101011010101",
		461 => "011000000101011010101",
		462 => "011010000100001010010",
		463 => "011010000100001010010",
		464 => "011010000100001010010",
		465 => "011000000101011010101",
		466 => "011000000101011010101",
		467 => "011000000101011010101",
		468 => "011001011101001010000",
		469 => "011001011101001010000",
		470 => "011001011101001010000",
		471 => "011000000101011010101",
		472 => "011000000101011010101",
		473 => "011000000101011010101",
		474 => "011010000100001010010",
		475 => "011010000100001010010",
		476 => "011010000100001010010",
		477 => "011000000101011010101",
		478 => "011000000101011010101",
		479 => "011000000101011010101",
		480 => "111011010100001010011",
		481 => "111011010100001010011",
		482 => "111011010100001010011",
		483 => "011000001101100010011",
		484 => "011000001101100010011",
		485 => "011000001101100010011",
		486 => "111011010100001010011",
		487 => "111011010100001010011",
		488 => "111011010100001010011",
		489 => "011000001101100010011",
		490 => "011000001101100010011",
		491 => "011000001101100010011",
		492 => "111011010100001010011",
		493 => "111011010100001010011",
		494 => "111011010100001010011",
		495 => "011000001101100010011",
		496 => "011000001101100010011",
		497 => "011000001101100010011",
		498 => "111011010100001010011",
		499 => "111011010100001010011",
		500 => "111011010100001010011",
		501 => "011000001101100010011",
		502 => "011000001101100010011",
		503 => "011000001101100010011",
		504 => "111011010100001010011",
		505 => "111011010100001010011",
		506 => "111011010100001010011",
		507 => "011000001101100010011",
		508 => "011000001101100010011",
		509 => "011000001101100010011",
		510 => "111011010100001010011",
		511 => "111011010100001010011",
		512 => "111011010100001010011",
		513 => "011000001101100010011",
		514 => "011000001101100010011",
		515 => "011000001101100010011",
		516 => "111011010100001010011",
		517 => "111011010100001010011",
		518 => "111011010100001010011",
		519 => "011000001101100010011",
		520 => "011000001101100010011",
		521 => "011000001101100010011",
		522 => "111011010100001010011",
		523 => "111011010100001010011",
		524 => "111011010100001010011",
		525 => "011000001101100010011",
		526 => "011000001101100010011",
		527 => "011000001101100010011",
		528 => "111011010100001010011",
		529 => "111011010100001010011",
		530 => "111011010100001010011",
		531 => "011000001101100010011",
		532 => "011000001101100010011",
		533 => "011000001101100010011",
		534 => "111011010100001010011",
		535 => "111011010100001010011",
		536 => "111011010100001010011",
		537 => "011000001101100010011",
		538 => "011000001101100010011",
		539 => "011000001101100010011",
		540 => "111011010100001010011",
		541 => "111011010100001010011",
		542 => "111011010100001010011",
		543 => "011000001101100010011",
		544 => "011000001101100010011",
		545 => "011000001101100010011",
		546 => "111011010100001010011",
		547 => "111011010100001010011",
		548 => "111011010100001010011",
		549 => "011000001101100010011",
		550 => "011000001101100010011",
		551 => "011000001101100010011",
		552 => "111011010100001010011",
		553 => "111011010100001010011",
		554 => "111011010100001010011",
		555 => "011000001101100010011",
		556 => "011000001101100010011",
		557 => "011000001101100010011",
		558 => "111011010100001010011",
		559 => "111011010100001010011",
		560 => "111011010100001010011",
		561 => "011000001101100010011",
		562 => "011000001101100010011",
		563 => "011000001101100010011",
		564 => "111011010100001010011",
		565 => "111011010100001010011",
		566 => "111011010100001010011",
		567 => "011000001101100010011",
		568 => "011000001101100010011",
		569 => "011000001101100010011",
		570 => "111011010100001010011",
		571 => "111011010100001010011",
		572 => "111011010100001010011",
		573 => "011000001101100010011",
		574 => "011000001101100010011",
		575 => "011000001101100010011",
		576 => "011011000100001110011",
		577 => "011011000100001110011",
		578 => "011011000100001110011",
		579 => "011011000100001110011",
		580 => "011011000100001110011",
		581 => "011011000100001110011",
		582 => "011011000100001110011",
		583 => "011011000100001110011",
		584 => "011011000100001110011",
		585 => "011011000100001110011",
		586 => "011011000100001110011",
		587 => "011011000100001110011",
		588 => "011011000100001110011",
		589 => "011011000100001110011",
		590 => "011011000100001110011",
		591 => "011011000100001110011",
		592 => "011011000100001110011",
		593 => "011011000100001110011",
		594 => "011011000100001110011",
		595 => "011011000100001110011",
		596 => "011011000100001110011",
		597 => "011011000100001110011",
		598 => "011011000100001110011",
		599 => "011011000100001110011",
		600 => "011011000100001110011",
		601 => "011011000100001110011",
		602 => "011011000100001110011",
		603 => "011011000100001110011",
		604 => "011011000100001110011",
		605 => "011011000100001110011",
		606 => "011011000100001110011",
		607 => "011011000100001110011",
		608 => "011011000100001110011",
		609 => "011011000100001110011",
		610 => "011011000100001110011",
		611 => "011011000100001110011",
		612 => "011011000100001110011",
		613 => "011011000100001110011",
		614 => "011011000100001110011",
		615 => "011011000100001110011",
		616 => "011011000100001110011",
		617 => "011011000100001110011",
		618 => "011011000100001110011",
		619 => "011011000100001110011",
		620 => "011011000100001110011",
		621 => "011011000100001110011",
		622 => "011011000100001110011",
		623 => "011011000100001110011",
		624 => "011011000100001110011",
		625 => "011011000100001110011",
		626 => "011011000100001110011",
		627 => "011011000100001110011",
		628 => "011011000100001110011",
		629 => "011011000100001110011",
		630 => "011011000100001110011",
		631 => "011011000100001110011",
		632 => "011011000100001110011",
		633 => "011011000100001110011",
		634 => "011011000100001110011",
		635 => "011011000100001110011",
		636 => "011011000100001110011",
		637 => "011011000100001110011",
		638 => "011011000100001110011",
		639 => "011011000100001110011",
		640 => "011011000100001110011",
		641 => "011011000100001110011",
		642 => "011011000100001110011",
		643 => "011011000100001110011",
		644 => "011011000100001110011",
		645 => "011011000100001110011",
		646 => "011011000100001110011",
		647 => "011011000100001110011",
		648 => "011011000100001110011",
		649 => "011011000100001110011",
		650 => "011011000100001110011",
		651 => "011011000100001110011",
		652 => "011011000100001110011",
		653 => "011011000100001110011",
		654 => "011011000100001110011",
		655 => "011011000100001110011",
		656 => "011011000100001110011",
		657 => "011011000100001110011",
		658 => "011011000100001110011",
		659 => "011011000100001110011",
		660 => "011011000100001110011",
		661 => "011011000100001110011",
		662 => "011011000100001110011",
		663 => "011011000100001110011",
		664 => "011011000100001110011",
		665 => "011011000100001110011",
		666 => "011011000100001110011",
		667 => "011011000100001110011",
		668 => "011011000100001110011",
		669 => "011011000100001110011",
		670 => "011011000100001110011",
		671 => "011011000100001110011",
		672 => "011000101100100010101",
		673 => "011000101100100010101",
		674 => "011000101100100010101",
		675 => "011000101100100010101",
		676 => "011000101100100010101",
		677 => "011000101100100010101",
		678 => "011000101100100010101",
		679 => "011000101100100010101",
		680 => "011000101100100010101",
		681 => "011000101100100010101",
		682 => "011000101100100010101",
		683 => "011000101100100010101",
		684 => "011000101100100010101",
		685 => "011000101100100010101",
		686 => "011000101100100010101",
		687 => "011000101100100010101",
		688 => "011000101100100010101",
		689 => "011000101100100010101",
		690 => "011000101100100010101",
		691 => "011000101100100010101",
		692 => "011000101100100010101",
		693 => "011000101100100010101",
		694 => "011000101100100010101",
		695 => "011000101100100010101",
		696 => "011000101100100010101",
		697 => "011000101100100010101",
		698 => "011000101100100010101",
		699 => "011000101100100010101",
		700 => "011000101100100010101",
		701 => "011000101100100010101",
		702 => "011000101100100010101",
		703 => "011000101100100010101",
		704 => "011000101100100010101",
		705 => "011000101100100010101",
		706 => "011000101100100010101",
		707 => "011000101100100010101",
		708 => "011000101100100010101",
		709 => "011000101100100010101",
		710 => "011000101100100010101",
		711 => "011000101100100010101",
		712 => "011000101100100010101",
		713 => "011000101100100010101",
		714 => "011000101100100010101",
		715 => "011000101100100010101",
		716 => "011000101100100010101",
		717 => "011000101100100010101",
		718 => "011000101100100010101",
		719 => "011000101100100010101",
		720 => "011000101100100010101",
		721 => "011000101100100010101",
		722 => "011000101100100010101",
		723 => "011000101100100010101",
		724 => "011000101100100010101",
		725 => "011000101100100010101",
		726 => "011000101100100010101",
		727 => "011000101100100010101",
		728 => "011000101100100010101",
		729 => "011000101100100010101",
		730 => "011000101100100010101",
		731 => "011000101100100010101",
		732 => "011000101100100010101",
		733 => "011000101100100010101",
		734 => "011000101100100010101",
		735 => "011000101100100010101",
		736 => "011000101100100010101",
		737 => "011000101100100010101",
		738 => "011000101100100010101",
		739 => "011000101100100010101",
		740 => "011000101100100010101",
		741 => "011000101100100010101",
		742 => "011000101100100010101",
		743 => "011000101100100010101",
		744 => "011000101100100010101",
		745 => "011000101100100010101",
		746 => "011000101100100010101",
		747 => "011000101100100010101",
		748 => "011000101100100010101",
		749 => "011000101100100010101",
		750 => "011000101100100010101",
		751 => "011000101100100010101",
		752 => "011000101100100010101",
		753 => "011000101100100010101",
		754 => "011000101100100010101",
		755 => "011000101100100010101",
		756 => "011000101100100010101",
		757 => "011000101100100010101",
		758 => "011000101100100010101",
		759 => "011000101100100010101",
		760 => "011000101100100010101",
		761 => "011000101100100010101",
		762 => "011000101100100010101",
		763 => "011000101100100010101",
		764 => "011000101100100010101",
		765 => "011000101100100010101",
		766 => "011000101100100010101",
		767 => "011000101100100010101",
		768 => "011000101100100110010",
		769 => "011000101100100110010",
		770 => "011000101100100110010",
		771 => "011000101100100110010",
		772 => "011000101100100110010",
		773 => "011000101100100110010",
		774 => "011000101100100110010",
		775 => "011000101100100110010",
		776 => "011000101100100110010",
		777 => "011000101100100110010",
		778 => "011000101100100110010",
		779 => "011000101100100110010",
		780 => "011000101100100110010",
		781 => "011000101100100110010",
		782 => "011000101100100110010",
		783 => "011000101100100110010",
		784 => "011000101100100110010",
		785 => "011000101100100110010",
		786 => "011000101100100110010",
		787 => "011000101100100110010",
		788 => "011000101100100110010",
		789 => "011000101100100110010",
		790 => "011000101100100110010",
		791 => "011000101100100110010",
		792 => "011000101100100110010",
		793 => "011000101100100110010",
		794 => "011000101100100110010",
		795 => "011000101100100110010",
		796 => "011000101100100110010",
		797 => "011000101100100110010",
		798 => "011000101100100110010",
		799 => "011000101100100110010",
		800 => "011000101100100110010",
		801 => "011000101100100110010",
		802 => "011000101100100110010",
		803 => "011000101100100110010",
		804 => "011000101100100110010",
		805 => "011000101100100110010",
		806 => "011000101100100110010",
		807 => "011000101100100110010",
		808 => "011000101100100110010",
		809 => "011000101100100110010",
		810 => "011000101100100110010",
		811 => "011000101100100110010",
		812 => "011000101100100110010",
		813 => "011000101100100110010",
		814 => "011000101100100110010",
		815 => "011000101100100110010",
		816 => "011000101100100110010",
		817 => "011000101100100110010",
		818 => "011000101100100110010",
		819 => "011000101100100110010",
		820 => "011000101100100110010",
		821 => "011000101100100110010",
		822 => "011000101100100110010",
		823 => "011000101100100110010",
		824 => "011000101100100110010",
		825 => "011000101100100110010",
		826 => "011000101100100110010",
		827 => "011000101100100110010",
		828 => "011000101100100110010",
		829 => "011000101100100110010",
		830 => "011000101100100110010",
		831 => "011000101100100110010",
		832 => "011000101100100110010",
		833 => "011000101100100110010",
		834 => "011000101100100110010",
		835 => "011000101100100110010",
		836 => "011000101100100110010",
		837 => "011000101100100110010",
		838 => "011000101100100110010",
		839 => "011000101100100110010",
		840 => "011000101100100110010",
		841 => "011000101100100110010",
		842 => "011000101100100110010",
		843 => "011000101100100110010",
		844 => "011000101100100110010",
		845 => "011000101100100110010",
		846 => "011000101100100110010",
		847 => "011000101100100110010",
		848 => "011000101100100110010",
		849 => "011000101100100110010",
		850 => "011000101100100110010",
		851 => "011000101100100110010",
		852 => "011000101100100110010",
		853 => "011000101100100110010",
		854 => "011000101100100110010",
		855 => "011000101100100110010",
		856 => "011000101100100110010",
		857 => "011000101100100110010",
		858 => "011000101100100110010",
		859 => "011000101100100110010",
		860 => "011000101100100110010",
		861 => "011000101100100110010",
		862 => "011000101100100110010",
		863 => "011000101100100110010");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;