library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT1 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT1;

architecture Behavioral of ROMFFT1 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 2 
	constant ROM_tb : ROM := (
		0 => "011100100111001110000",
		1 => "011100100111001110000",
		2 => "011100100111001110000",
		3 => "001011011101111010000",
		4 => "001011011101111010000",
		5 => "001011011101111010000",
		6 => "001000010100111010110",
		7 => "001000010100111010110",
		8 => "001000010100111010110",
		9 => "001010011100001010101",
		10 => "001010011100001010101",
		11 => "001010011100001010101",
		12 => "011000111100111010000",
		13 => "011000111100111010000",
		14 => "011000111100111010000",
		15 => "001001011100001010100",
		16 => "001001011100001010100",
		17 => "001001011100001010100",
		18 => "011000001100110010110",
		19 => "011000001100110010110",
		20 => "011000001100110010110",
		21 => "011000101100111110001",
		22 => "011000101100111110001",
		23 => "011000101100111110001",
		24 => "011000000100111010001",
		25 => "011000000100111010001",
		26 => "011000000100111010001",
		27 => "011000101100111010001",
		28 => "011000101100111010001",
		29 => "011000101100111010001",
		30 => "011000000100111010001",
		31 => "011000000100111010001",
		32 => "011000000100111010001",
		33 => "001000111100011110010",
		34 => "001000111100011110010",
		35 => "001000111100011110010",
		36 => "011000000100111010001",
		37 => "011000000100111010001",
		38 => "011000000100111010001",
		39 => "011000000101011010101",
		40 => "011000000101011010101",
		41 => "011000000101011010101",
		42 => "011000000101101010011",
		43 => "011000000101101010011",
		44 => "011000000101101010011",
		45 => "011000000110011010101",
		46 => "011000000110011010101",
		47 => "011000000110011010101",
		48 => "001000011110011011100",
		49 => "001000011110011011100",
		50 => "001000011110011011100",
		51 => "011011100100001110110",
		52 => "011011100100001110110",
		53 => "011011100100001110110",
		54 => "001000010100111010110",
		55 => "001000010100111010110",
		56 => "001000010100111010110",
		57 => "011010100100001010100",
		58 => "011010100100001010100",
		59 => "011010100100001010100",
		60 => "001000111100001010011",
		61 => "001000111100001010011",
		62 => "001000111100001010011",
		63 => "011010000100001010010",
		64 => "011010000100001010010",
		65 => "011010000100001010010",
		66 => "011000001100110010110",
		67 => "011000001100110010110",
		68 => "011000001100110010110",
		69 => "001000111100011110011",
		70 => "001000111100011110011",
		71 => "001000111100011110011",
		72 => "011000000100111010001",
		73 => "011000000100111010001",
		74 => "011000000100111010001",
		75 => "001000000100101110111",
		76 => "001000000100101110111",
		77 => "001000000100101110111",
		78 => "011000000100111010001",
		79 => "011000000100111010001",
		80 => "011000000100111010001",
		81 => "011001000100001010001",
		82 => "011001000100001010001",
		83 => "011001000100001010001",
		84 => "001000111100111010000",
		85 => "001000111100111010000",
		86 => "001000111100111010000",
		87 => "011000000101011010101",
		88 => "011000000101011010101",
		89 => "011000000101011010101",
		90 => "011011000100001110011",
		91 => "011011000100001110011",
		92 => "011011000100001110011",
		93 => "011000000110011010101",
		94 => "011000000110011010101",
		95 => "011000000110011010101",
		96 => "011011000110111010000",
		97 => "011011000110111010000",
		98 => "011011000110111010000",
		99 => "011010100100001110101",
		100 => "011010100100001110101",
		101 => "011010100100001110101",
		102 => "011001011100111010000",
		103 => "011001011100111010000",
		104 => "011001011100111010000",
		105 => "001000111100001110110",
		106 => "001000111100001110110",
		107 => "001000111100001110110",
		108 => "011001100100001110000",
		109 => "011001100100001110000",
		110 => "011001100100001110000",
		111 => "011000010100011010011",
		112 => "011000010100011010011",
		113 => "011000010100011010011",
		114 => "011000001100101010001",
		115 => "011000001100101010001",
		116 => "011000001100101010001",
		117 => "011000000101111010100",
		118 => "011000000101111010100",
		119 => "011000000101111010100",
		120 => "011101100101101110000",
		121 => "011101100101101110000",
		122 => "011101100101101110000",
		123 => "011010100100001110101",
		124 => "011010100100001110101",
		125 => "011010100100001110101",
		126 => "011001011100111010000",
		127 => "011001011100111010000",
		128 => "011001011100111010000",
		129 => "001000000101101010001",
		130 => "001000000101101010001",
		131 => "001000000101101010001",
		132 => "001000011100111010000",
		133 => "001000011100111010000",
		134 => "001000011100111010000",
		135 => "011000010100011010011",
		136 => "011000010100011010011",
		137 => "011000010100011010011",
		138 => "001000000100101110001",
		139 => "001000000100101110001",
		140 => "001000000100101110001",
		141 => "001010011101111010000",
		142 => "001010011101111010000",
		143 => "001010011101111010000",
		144 => "011011000110111010000",
		145 => "011011000110111010000",
		146 => "011011000110111010000",
		147 => "011010100100001110101",
		148 => "011010100100001110101",
		149 => "011010100100001110101",
		150 => "011001011100111010000",
		151 => "011001011100111010000",
		152 => "011001011100111010000",
		153 => "001000111100001110110",
		154 => "001000111100001110110",
		155 => "001000111100001110110",
		156 => "011001100100001110000",
		157 => "011001100100001110000",
		158 => "011001100100001110000",
		159 => "011000010100011010011",
		160 => "011000010100011010011",
		161 => "011000010100011010011",
		162 => "011000001100101010001",
		163 => "011000001100101010001",
		164 => "011000001100101010001",
		165 => "011000000101111010100",
		166 => "011000000101111010100",
		167 => "011000000101111010100",
		168 => "011101100101101110000",
		169 => "011101100101101110000",
		170 => "011101100101101110000",
		171 => "011010100100001110101",
		172 => "011010100100001110101",
		173 => "011010100100001110101",
		174 => "011001011100111010000",
		175 => "011001011100111010000",
		176 => "011001011100111010000",
		177 => "001000000101101010001",
		178 => "001000000101101010001",
		179 => "001000000101101010001",
		180 => "001000011100111010000",
		181 => "001000011100111010000",
		182 => "001000011100111010000",
		183 => "011000010100011010011",
		184 => "011000010100011010011",
		185 => "011000010100011010011",
		186 => "001000000100101110001",
		187 => "001000000100101110001",
		188 => "001000000100101110001",
		189 => "001010011101111010000",
		190 => "001010011101111010000",
		191 => "001010011101111010000",
		192 => "011000000110111110101",
		193 => "011000000110111110101",
		194 => "011000000110111110101",
		195 => "001000111100001110011",
		196 => "001000111100001110011",
		197 => "001000111100001110011",
		198 => "011001100100001110000",
		199 => "011001100100001110000",
		200 => "011001100100001110000",
		201 => "011010100100001110010",
		202 => "011010100100001110010",
		203 => "011010100100001110010",
		204 => "001010111100001011011",
		205 => "001010111100001011011",
		206 => "001010111100001011011",
		207 => "001000111100001110011",
		208 => "001000111100001110011",
		209 => "001000111100001110011",
		210 => "001000011100111010000",
		211 => "001000011100111010000",
		212 => "001000011100111010000",
		213 => "011000000101011010010",
		214 => "011000000101011010010",
		215 => "011000000101011010010",
		216 => "011000000110111110101",
		217 => "011000000110111110101",
		218 => "011000000110111110101",
		219 => "001000111100001110011",
		220 => "001000111100001110011",
		221 => "001000111100001110011",
		222 => "011001100100001110000",
		223 => "011001100100001110000",
		224 => "011001100100001110000",
		225 => "011010100100001110010",
		226 => "011010100100001110010",
		227 => "011010100100001110010",
		228 => "001010111100001011011",
		229 => "001010111100001011011",
		230 => "001010111100001011011",
		231 => "001000111100001110011",
		232 => "001000111100001110011",
		233 => "001000111100001110011",
		234 => "001000011100111010000",
		235 => "001000011100111010000",
		236 => "001000011100111010000",
		237 => "011000000101011010010",
		238 => "011000000101011010010",
		239 => "011000000101011010010",
		240 => "011000000110111110101",
		241 => "011000000110111110101",
		242 => "011000000110111110101",
		243 => "001000111100001110011",
		244 => "001000111100001110011",
		245 => "001000111100001110011",
		246 => "011001100100001110000",
		247 => "011001100100001110000",
		248 => "011001100100001110000",
		249 => "011010100100001110010",
		250 => "011010100100001110010",
		251 => "011010100100001110010",
		252 => "001010111100001011011",
		253 => "001010111100001011011",
		254 => "001010111100001011011",
		255 => "001000111100001110011",
		256 => "001000111100001110011",
		257 => "001000111100001110011",
		258 => "001000011100111010000",
		259 => "001000011100111010000",
		260 => "001000011100111010000",
		261 => "011000000101011010010",
		262 => "011000000101011010010",
		263 => "011000000101011010010",
		264 => "011000000110111110101",
		265 => "011000000110111110101",
		266 => "011000000110111110101",
		267 => "001000111100001110011",
		268 => "001000111100001110011",
		269 => "001000111100001110011",
		270 => "011001100100001110000",
		271 => "011001100100001110000",
		272 => "011001100100001110000",
		273 => "011010100100001110010",
		274 => "011010100100001110010",
		275 => "011010100100001110010",
		276 => "001010111100001011011",
		277 => "001010111100001011011",
		278 => "001010111100001011011",
		279 => "001000111100001110011",
		280 => "001000111100001110011",
		281 => "001000111100001110011",
		282 => "001000011100111010000",
		283 => "001000011100111010000",
		284 => "001000011100111010000",
		285 => "011000000101011010010",
		286 => "011000000101011010010",
		287 => "011000000101011010010",
		288 => "011000000110011110100",
		289 => "011000000110011110100",
		290 => "011000000110011110100",
		291 => "011001011100001010011",
		292 => "011001011100001010011",
		293 => "011001011100001010011",
		294 => "001010011100001011001",
		295 => "001010011100001011001",
		296 => "001010011100001011001",
		297 => "011001100100001110010",
		298 => "011001100100001110010",
		299 => "011001100100001110010",
		300 => "011000000110011110100",
		301 => "011000000110011110100",
		302 => "011000000110011110100",
		303 => "011001011100001010011",
		304 => "011001011100001010011",
		305 => "011001011100001010011",
		306 => "001010011100001011001",
		307 => "001010011100001011001",
		308 => "001010011100001011001",
		309 => "011001100100001110010",
		310 => "011001100100001110010",
		311 => "011001100100001110010",
		312 => "011000000110011110100",
		313 => "011000000110011110100",
		314 => "011000000110011110100",
		315 => "011001011100001010011",
		316 => "011001011100001010011",
		317 => "011001011100001010011",
		318 => "001010011100001011001",
		319 => "001010011100001011001",
		320 => "001010011100001011001",
		321 => "011001100100001110010",
		322 => "011001100100001110010",
		323 => "011001100100001110010",
		324 => "011000000110011110100",
		325 => "011000000110011110100",
		326 => "011000000110011110100",
		327 => "011001011100001010011",
		328 => "011001011100001010011",
		329 => "011001011100001010011",
		330 => "001010011100001011001",
		331 => "001010011100001011001",
		332 => "001010011100001011001",
		333 => "011001100100001110010",
		334 => "011001100100001110010",
		335 => "011001100100001110010",
		336 => "011000000110011110100",
		337 => "011000000110011110100",
		338 => "011000000110011110100",
		339 => "011001011100001010011",
		340 => "011001011100001010011",
		341 => "011001011100001010011",
		342 => "001010011100001011001",
		343 => "001010011100001011001",
		344 => "001010011100001011001",
		345 => "011001100100001110010",
		346 => "011001100100001110010",
		347 => "011001100100001110010",
		348 => "011000000110011110100",
		349 => "011000000110011110100",
		350 => "011000000110011110100",
		351 => "011001011100001010011",
		352 => "011001011100001010011",
		353 => "011001011100001010011",
		354 => "001010011100001011001",
		355 => "001010011100001011001",
		356 => "001010011100001011001",
		357 => "011001100100001110010",
		358 => "011001100100001110010",
		359 => "011001100100001110010",
		360 => "011000000110011110100",
		361 => "011000000110011110100",
		362 => "011000000110011110100",
		363 => "011001011100001010011",
		364 => "011001011100001010011",
		365 => "011001011100001010011",
		366 => "001010011100001011001",
		367 => "001010011100001011001",
		368 => "001010011100001011001",
		369 => "011001100100001110010",
		370 => "011001100100001110010",
		371 => "011001100100001110010",
		372 => "011000000110011110100",
		373 => "011000000110011110100",
		374 => "011000000110011110100",
		375 => "011001011100001010011",
		376 => "011001011100001010011",
		377 => "011001011100001010011",
		378 => "001010011100001011001",
		379 => "001010011100001011001",
		380 => "001010011100001011001",
		381 => "011001100100001110010",
		382 => "011001100100001110010",
		383 => "011001100100001110010",
		384 => "011000000101111110011",
		385 => "011000000101111110011",
		386 => "011000000101111110011",
		387 => "001001111100001010111",
		388 => "001001111100001010111",
		389 => "001001111100001010111",
		390 => "011000000101111110011",
		391 => "011000000101111110011",
		392 => "011000000101111110011",
		393 => "001001111100001010111",
		394 => "001001111100001010111",
		395 => "001001111100001010111",
		396 => "011000000101111110011",
		397 => "011000000101111110011",
		398 => "011000000101111110011",
		399 => "001001111100001010111",
		400 => "001001111100001010111",
		401 => "001001111100001010111",
		402 => "011000000101111110011",
		403 => "011000000101111110011",
		404 => "011000000101111110011",
		405 => "001001111100001010111",
		406 => "001001111100001010111",
		407 => "001001111100001010111",
		408 => "011000000101111110011",
		409 => "011000000101111110011",
		410 => "011000000101111110011",
		411 => "001001111100001010111",
		412 => "001001111100001010111",
		413 => "001001111100001010111",
		414 => "011000000101111110011",
		415 => "011000000101111110011",
		416 => "011000000101111110011",
		417 => "001001111100001010111",
		418 => "001001111100001010111",
		419 => "001001111100001010111",
		420 => "011000000101111110011",
		421 => "011000000101111110011",
		422 => "011000000101111110011",
		423 => "001001111100001010111",
		424 => "001001111100001010111",
		425 => "001001111100001010111",
		426 => "011000000101111110011",
		427 => "011000000101111110011",
		428 => "011000000101111110011",
		429 => "001001111100001010111",
		430 => "001001111100001010111",
		431 => "001001111100001010111",
		432 => "011000000101111110011",
		433 => "011000000101111110011",
		434 => "011000000101111110011",
		435 => "001001111100001010111",
		436 => "001001111100001010111",
		437 => "001001111100001010111",
		438 => "011000000101111110011",
		439 => "011000000101111110011",
		440 => "011000000101111110011",
		441 => "001001111100001010111",
		442 => "001001111100001010111",
		443 => "001001111100001010111",
		444 => "011000000101111110011",
		445 => "011000000101111110011",
		446 => "011000000101111110011",
		447 => "001001111100001010111",
		448 => "001001111100001010111",
		449 => "001001111100001010111",
		450 => "011000000101111110011",
		451 => "011000000101111110011",
		452 => "011000000101111110011",
		453 => "001001111100001010111",
		454 => "001001111100001010111",
		455 => "001001111100001010111",
		456 => "011000000101111110011",
		457 => "011000000101111110011",
		458 => "011000000101111110011",
		459 => "001001111100001010111",
		460 => "001001111100001010111",
		461 => "001001111100001010111",
		462 => "011000000101111110011",
		463 => "011000000101111110011",
		464 => "011000000101111110011",
		465 => "001001111100001010111",
		466 => "001001111100001010111",
		467 => "001001111100001010111",
		468 => "011000000101111110011",
		469 => "011000000101111110011",
		470 => "011000000101111110011",
		471 => "001001111100001010111",
		472 => "001001111100001010111",
		473 => "001001111100001010111",
		474 => "011000000101111110011",
		475 => "011000000101111110011",
		476 => "011000000101111110011",
		477 => "001001111100001010111",
		478 => "001001111100001010111",
		479 => "001001111100001010111",
		480 => "011010100100001110100",
		481 => "011010100100001110100",
		482 => "011010100100001110100",
		483 => "011010100100001110100",
		484 => "011010100100001110100",
		485 => "011010100100001110100",
		486 => "011010100100001110100",
		487 => "011010100100001110100",
		488 => "011010100100001110100",
		489 => "011010100100001110100",
		490 => "011010100100001110100",
		491 => "011010100100001110100",
		492 => "011010100100001110100",
		493 => "011010100100001110100",
		494 => "011010100100001110100",
		495 => "011010100100001110100",
		496 => "011010100100001110100",
		497 => "011010100100001110100",
		498 => "011010100100001110100",
		499 => "011010100100001110100",
		500 => "011010100100001110100",
		501 => "011010100100001110100",
		502 => "011010100100001110100",
		503 => "011010100100001110100",
		504 => "011010100100001110100",
		505 => "011010100100001110100",
		506 => "011010100100001110100",
		507 => "011010100100001110100",
		508 => "011010100100001110100",
		509 => "011010100100001110100",
		510 => "011010100100001110100",
		511 => "011010100100001110100",
		512 => "011010100100001110100",
		513 => "011010100100001110100",
		514 => "011010100100001110100",
		515 => "011010100100001110100",
		516 => "011010100100001110100",
		517 => "011010100100001110100",
		518 => "011010100100001110100",
		519 => "011010100100001110100",
		520 => "011010100100001110100",
		521 => "011010100100001110100",
		522 => "011010100100001110100",
		523 => "011010100100001110100",
		524 => "011010100100001110100",
		525 => "011010100100001110100",
		526 => "011010100100001110100",
		527 => "011010100100001110100",
		528 => "011010100100001110100",
		529 => "011010100100001110100",
		530 => "011010100100001110100",
		531 => "011010100100001110100",
		532 => "011010100100001110100",
		533 => "011010100100001110100",
		534 => "011010100100001110100",
		535 => "011010100100001110100",
		536 => "011010100100001110100",
		537 => "011010100100001110100",
		538 => "011010100100001110100",
		539 => "011010100100001110100",
		540 => "011010100100001110100",
		541 => "011010100100001110100",
		542 => "011010100100001110100",
		543 => "011010100100001110100",
		544 => "011010100100001110100",
		545 => "011010100100001110100",
		546 => "011010100100001110100",
		547 => "011010100100001110100",
		548 => "011010100100001110100",
		549 => "011010100100001110100",
		550 => "011010100100001110100",
		551 => "011010100100001110100",
		552 => "011010100100001110100",
		553 => "011010100100001110100",
		554 => "011010100100001110100",
		555 => "011010100100001110100",
		556 => "011010100100001110100",
		557 => "011010100100001110100",
		558 => "011010100100001110100",
		559 => "011010100100001110100",
		560 => "011010100100001110100",
		561 => "011010100100001110100",
		562 => "011010100100001110100",
		563 => "011010100100001110100",
		564 => "011010100100001110100",
		565 => "011010100100001110100",
		566 => "011010100100001110100",
		567 => "011010100100001110100",
		568 => "011010100100001110100",
		569 => "011010100100001110100",
		570 => "011010100100001110100",
		571 => "011010100100001110100",
		572 => "011010100100001110100",
		573 => "011010100100001110100",
		574 => "011010100100001110100",
		575 => "011010100100001110100",
		576 => "011001111100001010110",
		577 => "011001111100001010110",
		578 => "011001111100001010110",
		579 => "011001111100001010110",
		580 => "011001111100001010110",
		581 => "011001111100001010110",
		582 => "011001111100001010110",
		583 => "011001111100001010110",
		584 => "011001111100001010110",
		585 => "011001111100001010110",
		586 => "011001111100001010110",
		587 => "011001111100001010110",
		588 => "011001111100001010110",
		589 => "011001111100001010110",
		590 => "011001111100001010110",
		591 => "011001111100001010110",
		592 => "011001111100001010110",
		593 => "011001111100001010110",
		594 => "011001111100001010110",
		595 => "011001111100001010110",
		596 => "011001111100001010110",
		597 => "011001111100001010110",
		598 => "011001111100001010110",
		599 => "011001111100001010110",
		600 => "011001111100001010110",
		601 => "011001111100001010110",
		602 => "011001111100001010110",
		603 => "011001111100001010110",
		604 => "011001111100001010110",
		605 => "011001111100001010110",
		606 => "011001111100001010110",
		607 => "011001111100001010110",
		608 => "011001111100001010110",
		609 => "011001111100001010110",
		610 => "011001111100001010110",
		611 => "011001111100001010110",
		612 => "011001111100001010110",
		613 => "011001111100001010110",
		614 => "011001111100001010110",
		615 => "011001111100001010110",
		616 => "011001111100001010110",
		617 => "011001111100001010110",
		618 => "011001111100001010110",
		619 => "011001111100001010110",
		620 => "011001111100001010110",
		621 => "011001111100001010110",
		622 => "011001111100001010110",
		623 => "011001111100001010110",
		624 => "011001111100001010110",
		625 => "011001111100001010110",
		626 => "011001111100001010110",
		627 => "011001111100001010110",
		628 => "011001111100001010110",
		629 => "011001111100001010110",
		630 => "011001111100001010110",
		631 => "011001111100001010110",
		632 => "011001111100001010110",
		633 => "011001111100001010110",
		634 => "011001111100001010110",
		635 => "011001111100001010110",
		636 => "011001111100001010110",
		637 => "011001111100001010110",
		638 => "011001111100001010110",
		639 => "011001111100001010110",
		640 => "011001111100001010110",
		641 => "011001111100001010110",
		642 => "011001111100001010110",
		643 => "011001111100001010110",
		644 => "011001111100001010110",
		645 => "011001111100001010110",
		646 => "011001111100001010110",
		647 => "011001111100001010110",
		648 => "011001111100001010110",
		649 => "011001111100001010110",
		650 => "011001111100001010110",
		651 => "011001111100001010110",
		652 => "011001111100001010110",
		653 => "011001111100001010110",
		654 => "011001111100001010110",
		655 => "011001111100001010110",
		656 => "011001111100001010110",
		657 => "011001111100001010110",
		658 => "011001111100001010110",
		659 => "011001111100001010110",
		660 => "011001111100001010110",
		661 => "011001111100001010110",
		662 => "011001111100001010110",
		663 => "011001111100001010110",
		664 => "011001111100001010110",
		665 => "011001111100001010110",
		666 => "011001111100001010110",
		667 => "011001111100001010110",
		668 => "011001111100001010110",
		669 => "011001111100001010110",
		670 => "011001111100001010110",
		671 => "011001111100001010110",
		672 => "011000101100100010101",
		673 => "011000101100100010101",
		674 => "011000101100100010101",
		675 => "011000101100100010101",
		676 => "011000101100100010101",
		677 => "011000101100100010101",
		678 => "011000101100100010101",
		679 => "011000101100100010101",
		680 => "011000101100100010101",
		681 => "011000101100100010101",
		682 => "011000101100100010101",
		683 => "011000101100100010101",
		684 => "011000101100100010101",
		685 => "011000101100100010101",
		686 => "011000101100100010101",
		687 => "011000101100100010101",
		688 => "011000101100100010101",
		689 => "011000101100100010101",
		690 => "011000101100100010101",
		691 => "011000101100100010101",
		692 => "011000101100100010101",
		693 => "011000101100100010101",
		694 => "011000101100100010101",
		695 => "011000101100100010101",
		696 => "011000101100100010101",
		697 => "011000101100100010101",
		698 => "011000101100100010101",
		699 => "011000101100100010101",
		700 => "011000101100100010101",
		701 => "011000101100100010101",
		702 => "011000101100100010101",
		703 => "011000101100100010101",
		704 => "011000101100100010101",
		705 => "011000101100100010101",
		706 => "011000101100100010101",
		707 => "011000101100100010101",
		708 => "011000101100100010101",
		709 => "011000101100100010101",
		710 => "011000101100100010101",
		711 => "011000101100100010101",
		712 => "011000101100100010101",
		713 => "011000101100100010101",
		714 => "011000101100100010101",
		715 => "011000101100100010101",
		716 => "011000101100100010101",
		717 => "011000101100100010101",
		718 => "011000101100100010101",
		719 => "011000101100100010101",
		720 => "011000101100100010101",
		721 => "011000101100100010101",
		722 => "011000101100100010101",
		723 => "011000101100100010101",
		724 => "011000101100100010101",
		725 => "011000101100100010101",
		726 => "011000101100100010101",
		727 => "011000101100100010101",
		728 => "011000101100100010101",
		729 => "011000101100100010101",
		730 => "011000101100100010101",
		731 => "011000101100100010101",
		732 => "011000101100100010101",
		733 => "011000101100100010101",
		734 => "011000101100100010101",
		735 => "011000101100100010101",
		736 => "011000101100100010101",
		737 => "011000101100100010101",
		738 => "011000101100100010101",
		739 => "011000101100100010101",
		740 => "011000101100100010101",
		741 => "011000101100100010101",
		742 => "011000101100100010101",
		743 => "011000101100100010101",
		744 => "011000101100100010101",
		745 => "011000101100100010101",
		746 => "011000101100100010101",
		747 => "011000101100100010101",
		748 => "011000101100100010101",
		749 => "011000101100100010101",
		750 => "011000101100100010101",
		751 => "011000101100100010101",
		752 => "011000101100100010101",
		753 => "011000101100100010101",
		754 => "011000101100100010101",
		755 => "011000101100100010101",
		756 => "011000101100100010101",
		757 => "011000101100100010101",
		758 => "011000101100100010101",
		759 => "011000101100100010101",
		760 => "011000101100100010101",
		761 => "011000101100100010101",
		762 => "011000101100100010101",
		763 => "011000101100100010101",
		764 => "011000101100100010101",
		765 => "011000101100100010101",
		766 => "011000101100100010101",
		767 => "011000101100100010101",
		768 => "011000101100100110010",
		769 => "011000101100100110010",
		770 => "011000101100100110010",
		771 => "011000101100100110010",
		772 => "011000101100100110010",
		773 => "011000101100100110010",
		774 => "011000101100100110010",
		775 => "011000101100100110010",
		776 => "011000101100100110010",
		777 => "011000101100100110010",
		778 => "011000101100100110010",
		779 => "011000101100100110010",
		780 => "011000101100100110010",
		781 => "011000101100100110010",
		782 => "011000101100100110010",
		783 => "011000101100100110010",
		784 => "011000101100100110010",
		785 => "011000101100100110010",
		786 => "011000101100100110010",
		787 => "011000101100100110010",
		788 => "011000101100100110010",
		789 => "011000101100100110010",
		790 => "011000101100100110010",
		791 => "011000101100100110010",
		792 => "011000101100100110010",
		793 => "011000101100100110010",
		794 => "011000101100100110010",
		795 => "011000101100100110010",
		796 => "011000101100100110010",
		797 => "011000101100100110010",
		798 => "011000101100100110010",
		799 => "011000101100100110010",
		800 => "011000101100100110010",
		801 => "011000101100100110010",
		802 => "011000101100100110010",
		803 => "011000101100100110010",
		804 => "011000101100100110010",
		805 => "011000101100100110010",
		806 => "011000101100100110010",
		807 => "011000101100100110010",
		808 => "011000101100100110010",
		809 => "011000101100100110010",
		810 => "011000101100100110010",
		811 => "011000101100100110010",
		812 => "011000101100100110010",
		813 => "011000101100100110010",
		814 => "011000101100100110010",
		815 => "011000101100100110010",
		816 => "011000101100100110010",
		817 => "011000101100100110010",
		818 => "011000101100100110010",
		819 => "011000101100100110010",
		820 => "011000101100100110010",
		821 => "011000101100100110010",
		822 => "011000101100100110010",
		823 => "011000101100100110010",
		824 => "011000101100100110010",
		825 => "011000101100100110010",
		826 => "011000101100100110010",
		827 => "011000101100100110010",
		828 => "011000101100100110010",
		829 => "011000101100100110010",
		830 => "011000101100100110010",
		831 => "011000101100100110010",
		832 => "011000101100100110010",
		833 => "011000101100100110010",
		834 => "011000101100100110010",
		835 => "011000101100100110010",
		836 => "011000101100100110010",
		837 => "011000101100100110010",
		838 => "011000101100100110010",
		839 => "011000101100100110010",
		840 => "011000101100100110010",
		841 => "011000101100100110010",
		842 => "011000101100100110010",
		843 => "011000101100100110010",
		844 => "011000101100100110010",
		845 => "011000101100100110010",
		846 => "011000101100100110010",
		847 => "011000101100100110010",
		848 => "011000101100100110010",
		849 => "011000101100100110010",
		850 => "011000101100100110010",
		851 => "011000101100100110010",
		852 => "011000101100100110010",
		853 => "011000101100100110010",
		854 => "011000101100100110010",
		855 => "011000101100100110010",
		856 => "011000101100100110010",
		857 => "011000101100100110010",
		858 => "011000101100100110010",
		859 => "011000101100100110010",
		860 => "011000101100100110010",
		861 => "011000101100100110010",
		862 => "011000101100100110010",
		863 => "011000101100100110010");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;