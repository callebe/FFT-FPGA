library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT15 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT15;

architecture Behavioral of ROMFFT15 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 16 
	constant ROM_tb : ROM := (
		0 => "001010111100001011001",
		1 => "001010111100001011001",
		2 => "001010111100001011001",
		3 => "001001111100001010110",
		4 => "001001111100001010110",
		5 => "001001111100001010110",
		6 => "001010111100001010101",
		7 => "001010111100001010101",
		8 => "001010111100001010101",
		9 => "011000000100111110001",
		10 => "011000000100111110001",
		11 => "011000000100111110001",
		12 => "011000101100101010001",
		13 => "011000101100101010001",
		14 => "011000101100101010001",
		15 => "001000111100001010011",
		16 => "001000111100001010011",
		17 => "001000111100001010011",
		18 => "001000111100011110011",
		19 => "001000111100011110011",
		20 => "001000111100011110011",
		21 => "001000111100001010011",
		22 => "001000111100001010011",
		23 => "001000111100001010011",
		24 => "011000101100111010001",
		25 => "011000101100111010001",
		26 => "011000101100111010001",
		27 => "011000001100110010110",
		28 => "011000001100110010110",
		29 => "011000001100110010110",
		30 => "011000000101001010010",
		31 => "011000000101001010010",
		32 => "011000000101001010010",
		33 => "011001100100001110001",
		34 => "011001100100001110001",
		35 => "011001100100001110001",
		36 => "011000000101011010100",
		37 => "011000000101011010100",
		38 => "011000000101011010100",
		39 => "011000010100111010110",
		40 => "011000010100111010110",
		41 => "011000010100111010110",
		42 => "001011011100001010111",
		43 => "001011011100001010111",
		44 => "001011011100001010111",
		45 => "011100100111001010000",
		46 => "011100100111001010000",
		47 => "011100100111001010000",
		48 => "011100100100001010101",
		49 => "011100100100001010101",
		50 => "011100100100001010101",
		51 => "011011000100001010011",
		52 => "011011000100001010011",
		53 => "011011000100001010011",
		54 => "011010100100001010101",
		55 => "011010100100001010101",
		56 => "011010100100001010101",
		57 => "001000111100001010011",
		58 => "001000111100001010011",
		59 => "001000111100001010011",
		60 => "011001000100001110001",
		61 => "011001000100001110001",
		62 => "011001000100001110001",
		63 => "011001100100001010001",
		64 => "011001100100001010001",
		65 => "011001100100001010001",
		66 => "001000100100111010001",
		67 => "001000100100111010001",
		68 => "001000100100111010001",
		69 => "011010100100001010010",
		70 => "011010100100001010010",
		71 => "011010100100001010010",
		72 => "011000101100111010001",
		73 => "011000101100111010001",
		74 => "011000101100111010001",
		75 => "011000001100110010110",
		76 => "011000001100110010110",
		77 => "011000001100110010110",
		78 => "011010000100001110010",
		79 => "011010000100001110010",
		80 => "011010000100001110010",
		81 => "001000111100111010000",
		82 => "001000111100111010000",
		83 => "001000111100111010000",
		84 => "011000000101011010100",
		85 => "011000000101011010100",
		86 => "011000000101011010100",
		87 => "011000010100111010110",
		88 => "011000010100111010110",
		89 => "011000010100111010110",
		90 => "011011100100001010110",
		91 => "011011100100001010110",
		92 => "011011100100001010110",
		93 => "001000011111001011001",
		94 => "001000011111001011001",
		95 => "001000011111001011001",
		96 => "001010011100001010111",
		97 => "001010011100001010111",
		98 => "001010011100001010111",
		99 => "011000110100001010010",
		100 => "011000110100001010010",
		101 => "011000110100001010010",
		102 => "001000100100111110000",
		103 => "001000100100111110000",
		104 => "001000100100111110000",
		105 => "011000011100111010000",
		106 => "011000011100111010000",
		107 => "011000011100111010000",
		108 => "011001111100001010011",
		109 => "011001111100001010011",
		110 => "011001111100001010011",
		111 => "011001100100001110010",
		112 => "011001100100001110010",
		113 => "011001100100001110010",
		114 => "001010111100001010101",
		115 => "001010111100001010101",
		116 => "001010111100001010101",
		117 => "001000011101101011011",
		118 => "001000011101101011011",
		119 => "001000011101101011011",
		120 => "011011100100001010100",
		121 => "011011100100001010100",
		122 => "011011100100001010100",
		123 => "001000111100001110010",
		124 => "001000111100001110010",
		125 => "001000111100001110010",
		126 => "001000010100011010011",
		127 => "001000010100011010011",
		128 => "001000010100011010011",
		129 => "011001000100001110100",
		130 => "011001000100001110100",
		131 => "011001000100001110100",
		132 => "011001100100001110011",
		133 => "011001100100001110011",
		134 => "011001100100001110011",
		135 => "011000000100111010010",
		136 => "011000000100111010010",
		137 => "011000000100111010010",
		138 => "011010100100001010101",
		139 => "011010100100001010101",
		140 => "011010100100001010101",
		141 => "011101100101101010000",
		142 => "011101100101101010000",
		143 => "011101100101101010000",
		144 => "001010011100001010111",
		145 => "001010011100001010111",
		146 => "001010011100001010111",
		147 => "011000110100001010010",
		148 => "011000110100001010010",
		149 => "011000110100001010010",
		150 => "001000100100111110000",
		151 => "001000100100111110000",
		152 => "001000100100111110000",
		153 => "011000011100111010000",
		154 => "011000011100111010000",
		155 => "011000011100111010000",
		156 => "011001111100001010011",
		157 => "011001111100001010011",
		158 => "011001111100001010011",
		159 => "011001100100001110010",
		160 => "011001100100001110010",
		161 => "011001100100001110010",
		162 => "001010111100001010101",
		163 => "001010111100001010101",
		164 => "001010111100001010101",
		165 => "001000011101101011011",
		166 => "001000011101101011011",
		167 => "001000011101101011011",
		168 => "011011100100001010100",
		169 => "011011100100001010100",
		170 => "011011100100001010100",
		171 => "001000111100001110010",
		172 => "001000111100001110010",
		173 => "001000111100001110010",
		174 => "001000010100011010011",
		175 => "001000010100011010011",
		176 => "001000010100011010011",
		177 => "011001000100001110100",
		178 => "011001000100001110100",
		179 => "011001000100001110100",
		180 => "011001100100001110011",
		181 => "011001100100001110011",
		182 => "011001100100001110011",
		183 => "011000000100111010010",
		184 => "011000000100111010010",
		185 => "011000000100111010010",
		186 => "011010100100001010101",
		187 => "011010100100001010101",
		188 => "011010100100001010101",
		189 => "011101100101101010000",
		190 => "011101100101101010000",
		191 => "011101100101101010000",
		192 => "011010100100001010010",
		193 => "011010100100001010010",
		194 => "011010100100001010010",
		195 => "011000011100111010000",
		196 => "011000011100111010000",
		197 => "011000011100111010000",
		198 => "001000110100001010011",
		199 => "001000110100001010011",
		200 => "001000110100001010011",
		201 => "011000000110111010101",
		202 => "011000000110111010101",
		203 => "011000000110111010101",
		204 => "011010100100001010010",
		205 => "011010100100001010010",
		206 => "011010100100001010010",
		207 => "011001000100001110100",
		208 => "011001000100001110100",
		209 => "011001000100001110100",
		210 => "011000101100100110100",
		211 => "011000101100100110100",
		212 => "011000101100100110100",
		213 => "001000011110101010111",
		214 => "001000011110101010111",
		215 => "001000011110101010111",
		216 => "011010100100001010010",
		217 => "011010100100001010010",
		218 => "011010100100001010010",
		219 => "011000011100111010000",
		220 => "011000011100111010000",
		221 => "011000011100111010000",
		222 => "001000110100001010011",
		223 => "001000110100001010011",
		224 => "001000110100001010011",
		225 => "011000000110111010101",
		226 => "011000000110111010101",
		227 => "011000000110111010101",
		228 => "011010100100001010010",
		229 => "011010100100001010010",
		230 => "011010100100001010010",
		231 => "011001000100001110100",
		232 => "011001000100001110100",
		233 => "011001000100001110100",
		234 => "011000101100100110100",
		235 => "011000101100100110100",
		236 => "011000101100100110100",
		237 => "001000011110101010111",
		238 => "001000011110101010111",
		239 => "001000011110101010111",
		240 => "011010100100001010010",
		241 => "011010100100001010010",
		242 => "011010100100001010010",
		243 => "011000011100111010000",
		244 => "011000011100111010000",
		245 => "011000011100111010000",
		246 => "001000110100001010011",
		247 => "001000110100001010011",
		248 => "001000110100001010011",
		249 => "011000000110111010101",
		250 => "011000000110111010101",
		251 => "011000000110111010101",
		252 => "011010100100001010010",
		253 => "011010100100001010010",
		254 => "011010100100001010010",
		255 => "011001000100001110100",
		256 => "011001000100001110100",
		257 => "011001000100001110100",
		258 => "011000101100100110100",
		259 => "011000101100100110100",
		260 => "011000101100100110100",
		261 => "001000011110101010111",
		262 => "001000011110101010111",
		263 => "001000011110101010111",
		264 => "011010100100001010010",
		265 => "011010100100001010010",
		266 => "011010100100001010010",
		267 => "011000011100111010000",
		268 => "011000011100111010000",
		269 => "011000011100111010000",
		270 => "001000110100001010011",
		271 => "001000110100001010011",
		272 => "001000110100001010011",
		273 => "011000000110111010101",
		274 => "011000000110111010101",
		275 => "011000000110111010101",
		276 => "011010100100001010010",
		277 => "011010100100001010010",
		278 => "011010100100001010010",
		279 => "011001000100001110100",
		280 => "011001000100001110100",
		281 => "011001000100001110100",
		282 => "011000101100100110100",
		283 => "011000101100100110100",
		284 => "011000101100100110100",
		285 => "001000011110101010111",
		286 => "001000011110101010111",
		287 => "001000011110101010111",
		288 => "011001011100111010000",
		289 => "011001011100111010000",
		290 => "011001011100111010000",
		291 => "011000000110011010100",
		292 => "011000000110011010100",
		293 => "011000000110011010100",
		294 => "011001100100001010010",
		295 => "011001100100001010010",
		296 => "011001100100001010010",
		297 => "001010011110011010000",
		298 => "001010011110011010000",
		299 => "001010011110011010000",
		300 => "011001011100111010000",
		301 => "011001011100111010000",
		302 => "011001011100111010000",
		303 => "011000000110011010100",
		304 => "011000000110011010100",
		305 => "011000000110011010100",
		306 => "011001100100001010010",
		307 => "011001100100001010010",
		308 => "011001100100001010010",
		309 => "001010011110011010000",
		310 => "001010011110011010000",
		311 => "001010011110011010000",
		312 => "011001011100111010000",
		313 => "011001011100111010000",
		314 => "011001011100111010000",
		315 => "011000000110011010100",
		316 => "011000000110011010100",
		317 => "011000000110011010100",
		318 => "011001100100001010010",
		319 => "011001100100001010010",
		320 => "011001100100001010010",
		321 => "001010011110011010000",
		322 => "001010011110011010000",
		323 => "001010011110011010000",
		324 => "011001011100111010000",
		325 => "011001011100111010000",
		326 => "011001011100111010000",
		327 => "011000000110011010100",
		328 => "011000000110011010100",
		329 => "011000000110011010100",
		330 => "011001100100001010010",
		331 => "011001100100001010010",
		332 => "011001100100001010010",
		333 => "001010011110011010000",
		334 => "001010011110011010000",
		335 => "001010011110011010000",
		336 => "011001011100111010000",
		337 => "011001011100111010000",
		338 => "011001011100111010000",
		339 => "011000000110011010100",
		340 => "011000000110011010100",
		341 => "011000000110011010100",
		342 => "011001100100001010010",
		343 => "011001100100001010010",
		344 => "011001100100001010010",
		345 => "001010011110011010000",
		346 => "001010011110011010000",
		347 => "001010011110011010000",
		348 => "011001011100111010000",
		349 => "011001011100111010000",
		350 => "011001011100111010000",
		351 => "011000000110011010100",
		352 => "011000000110011010100",
		353 => "011000000110011010100",
		354 => "011001100100001010010",
		355 => "011001100100001010010",
		356 => "011001100100001010010",
		357 => "001010011110011010000",
		358 => "001010011110011010000",
		359 => "001010011110011010000",
		360 => "011001011100111010000",
		361 => "011001011100111010000",
		362 => "011001011100111010000",
		363 => "011000000110011010100",
		364 => "011000000110011010100",
		365 => "011000000110011010100",
		366 => "011001100100001010010",
		367 => "011001100100001010010",
		368 => "011001100100001010010",
		369 => "001010011110011010000",
		370 => "001010011110011010000",
		371 => "001010011110011010000",
		372 => "011001011100111010000",
		373 => "011001011100111010000",
		374 => "011001011100111010000",
		375 => "011000000110011010100",
		376 => "011000000110011010100",
		377 => "011000000110011010100",
		378 => "011001100100001010010",
		379 => "011001100100001010010",
		380 => "011001100100001010010",
		381 => "001010011110011010000",
		382 => "001010011110011010000",
		383 => "001010011110011010000",
		384 => "011011100100001110011",
		385 => "011011100100001110011",
		386 => "011011100100001110011",
		387 => "011000000101111010011",
		388 => "011000000101111010011",
		389 => "011000000101111010011",
		390 => "011011100100001110011",
		391 => "011011100100001110011",
		392 => "011011100100001110011",
		393 => "011000000101111010011",
		394 => "011000000101111010011",
		395 => "011000000101111010011",
		396 => "011011100100001110011",
		397 => "011011100100001110011",
		398 => "011011100100001110011",
		399 => "011000000101111010011",
		400 => "011000000101111010011",
		401 => "011000000101111010011",
		402 => "011011100100001110011",
		403 => "011011100100001110011",
		404 => "011011100100001110011",
		405 => "011000000101111010011",
		406 => "011000000101111010011",
		407 => "011000000101111010011",
		408 => "011011100100001110011",
		409 => "011011100100001110011",
		410 => "011011100100001110011",
		411 => "011000000101111010011",
		412 => "011000000101111010011",
		413 => "011000000101111010011",
		414 => "011011100100001110011",
		415 => "011011100100001110011",
		416 => "011011100100001110011",
		417 => "011000000101111010011",
		418 => "011000000101111010011",
		419 => "011000000101111010011",
		420 => "011011100100001110011",
		421 => "011011100100001110011",
		422 => "011011100100001110011",
		423 => "011000000101111010011",
		424 => "011000000101111010011",
		425 => "011000000101111010011",
		426 => "011011100100001110011",
		427 => "011011100100001110011",
		428 => "011011100100001110011",
		429 => "011000000101111010011",
		430 => "011000000101111010011",
		431 => "011000000101111010011",
		432 => "011011100100001110011",
		433 => "011011100100001110011",
		434 => "011011100100001110011",
		435 => "011000000101111010011",
		436 => "011000000101111010011",
		437 => "011000000101111010011",
		438 => "011011100100001110011",
		439 => "011011100100001110011",
		440 => "011011100100001110011",
		441 => "011000000101111010011",
		442 => "011000000101111010011",
		443 => "011000000101111010011",
		444 => "011011100100001110011",
		445 => "011011100100001110011",
		446 => "011011100100001110011",
		447 => "011000000101111010011",
		448 => "011000000101111010011",
		449 => "011000000101111010011",
		450 => "011011100100001110011",
		451 => "011011100100001110011",
		452 => "011011100100001110011",
		453 => "011000000101111010011",
		454 => "011000000101111010011",
		455 => "011000000101111010011",
		456 => "011011100100001110011",
		457 => "011011100100001110011",
		458 => "011011100100001110011",
		459 => "011000000101111010011",
		460 => "011000000101111010011",
		461 => "011000000101111010011",
		462 => "011011100100001110011",
		463 => "011011100100001110011",
		464 => "011011100100001110011",
		465 => "011000000101111010011",
		466 => "011000000101111010011",
		467 => "011000000101111010011",
		468 => "011011100100001110011",
		469 => "011011100100001110011",
		470 => "011011100100001110011",
		471 => "011000000101111010011",
		472 => "011000000101111010011",
		473 => "011000000101111010011",
		474 => "011011100100001110011",
		475 => "011011100100001110011",
		476 => "011011100100001110011",
		477 => "011000000101111010011",
		478 => "011000000101111010011",
		479 => "011000000101111010011",
		480 => "011010100100001010100",
		481 => "011010100100001010100",
		482 => "011010100100001010100",
		483 => "011010100100001010100",
		484 => "011010100100001010100",
		485 => "011010100100001010100",
		486 => "011010100100001010100",
		487 => "011010100100001010100",
		488 => "011010100100001010100",
		489 => "011010100100001010100",
		490 => "011010100100001010100",
		491 => "011010100100001010100",
		492 => "011010100100001010100",
		493 => "011010100100001010100",
		494 => "011010100100001010100",
		495 => "011010100100001010100",
		496 => "011010100100001010100",
		497 => "011010100100001010100",
		498 => "011010100100001010100",
		499 => "011010100100001010100",
		500 => "011010100100001010100",
		501 => "011010100100001010100",
		502 => "011010100100001010100",
		503 => "011010100100001010100",
		504 => "011010100100001010100",
		505 => "011010100100001010100",
		506 => "011010100100001010100",
		507 => "011010100100001010100",
		508 => "011010100100001010100",
		509 => "011010100100001010100",
		510 => "011010100100001010100",
		511 => "011010100100001010100",
		512 => "011010100100001010100",
		513 => "011010100100001010100",
		514 => "011010100100001010100",
		515 => "011010100100001010100",
		516 => "011010100100001010100",
		517 => "011010100100001010100",
		518 => "011010100100001010100",
		519 => "011010100100001010100",
		520 => "011010100100001010100",
		521 => "011010100100001010100",
		522 => "011010100100001010100",
		523 => "011010100100001010100",
		524 => "011010100100001010100",
		525 => "011010100100001010100",
		526 => "011010100100001010100",
		527 => "011010100100001010100",
		528 => "011010100100001010100",
		529 => "011010100100001010100",
		530 => "011010100100001010100",
		531 => "011010100100001010100",
		532 => "011010100100001010100",
		533 => "011010100100001010100",
		534 => "011010100100001010100",
		535 => "011010100100001010100",
		536 => "011010100100001010100",
		537 => "011010100100001010100",
		538 => "011010100100001010100",
		539 => "011010100100001010100",
		540 => "011010100100001010100",
		541 => "011010100100001010100",
		542 => "011010100100001010100",
		543 => "011010100100001010100",
		544 => "011010100100001010100",
		545 => "011010100100001010100",
		546 => "011010100100001010100",
		547 => "011010100100001010100",
		548 => "011010100100001010100",
		549 => "011010100100001010100",
		550 => "011010100100001010100",
		551 => "011010100100001010100",
		552 => "011010100100001010100",
		553 => "011010100100001010100",
		554 => "011010100100001010100",
		555 => "011010100100001010100",
		556 => "011010100100001010100",
		557 => "011010100100001010100",
		558 => "011010100100001010100",
		559 => "011010100100001010100",
		560 => "011010100100001010100",
		561 => "011010100100001010100",
		562 => "011010100100001010100",
		563 => "011010100100001010100",
		564 => "011010100100001010100",
		565 => "011010100100001010100",
		566 => "011010100100001010100",
		567 => "011010100100001010100",
		568 => "011010100100001010100",
		569 => "011010100100001010100",
		570 => "011010100100001010100",
		571 => "011010100100001010100",
		572 => "011010100100001010100",
		573 => "011010100100001010100",
		574 => "011010100100001010100",
		575 => "011010100100001010100",
		576 => "001000111100111010000",
		577 => "001000111100111010000",
		578 => "001000111100111010000",
		579 => "001000111100111010000",
		580 => "001000111100111010000",
		581 => "001000111100111010000",
		582 => "001000111100111010000",
		583 => "001000111100111010000",
		584 => "001000111100111010000",
		585 => "001000111100111010000",
		586 => "001000111100111010000",
		587 => "001000111100111010000",
		588 => "001000111100111010000",
		589 => "001000111100111010000",
		590 => "001000111100111010000",
		591 => "001000111100111010000",
		592 => "001000111100111010000",
		593 => "001000111100111010000",
		594 => "001000111100111010000",
		595 => "001000111100111010000",
		596 => "001000111100111010000",
		597 => "001000111100111010000",
		598 => "001000111100111010000",
		599 => "001000111100111010000",
		600 => "001000111100111010000",
		601 => "001000111100111010000",
		602 => "001000111100111010000",
		603 => "001000111100111010000",
		604 => "001000111100111010000",
		605 => "001000111100111010000",
		606 => "001000111100111010000",
		607 => "001000111100111010000",
		608 => "001000111100111010000",
		609 => "001000111100111010000",
		610 => "001000111100111010000",
		611 => "001000111100111010000",
		612 => "001000111100111010000",
		613 => "001000111100111010000",
		614 => "001000111100111010000",
		615 => "001000111100111010000",
		616 => "001000111100111010000",
		617 => "001000111100111010000",
		618 => "001000111100111010000",
		619 => "001000111100111010000",
		620 => "001000111100111010000",
		621 => "001000111100111010000",
		622 => "001000111100111010000",
		623 => "001000111100111010000",
		624 => "001000111100111010000",
		625 => "001000111100111010000",
		626 => "001000111100111010000",
		627 => "001000111100111010000",
		628 => "001000111100111010000",
		629 => "001000111100111010000",
		630 => "001000111100111010000",
		631 => "001000111100111010000",
		632 => "001000111100111010000",
		633 => "001000111100111010000",
		634 => "001000111100111010000",
		635 => "001000111100111010000",
		636 => "001000111100111010000",
		637 => "001000111100111010000",
		638 => "001000111100111010000",
		639 => "001000111100111010000",
		640 => "001000111100111010000",
		641 => "001000111100111010000",
		642 => "001000111100111010000",
		643 => "001000111100111010000",
		644 => "001000111100111010000",
		645 => "001000111100111010000",
		646 => "001000111100111010000",
		647 => "001000111100111010000",
		648 => "001000111100111010000",
		649 => "001000111100111010000",
		650 => "001000111100111010000",
		651 => "001000111100111010000",
		652 => "001000111100111010000",
		653 => "001000111100111010000",
		654 => "001000111100111010000",
		655 => "001000111100111010000",
		656 => "001000111100111010000",
		657 => "001000111100111010000",
		658 => "001000111100111010000",
		659 => "001000111100111010000",
		660 => "001000111100111010000",
		661 => "001000111100111010000",
		662 => "001000111100111010000",
		663 => "001000111100111010000",
		664 => "001000111100111010000",
		665 => "001000111100111010000",
		666 => "001000111100111010000",
		667 => "001000111100111010000",
		668 => "001000111100111010000",
		669 => "001000111100111010000",
		670 => "001000111100111010000",
		671 => "001000111100111010000",
		672 => "011000101100100010101",
		673 => "011000101100100010101",
		674 => "011000101100100010101",
		675 => "011000101100100010101",
		676 => "011000101100100010101",
		677 => "011000101100100010101",
		678 => "011000101100100010101",
		679 => "011000101100100010101",
		680 => "011000101100100010101",
		681 => "011000101100100010101",
		682 => "011000101100100010101",
		683 => "011000101100100010101",
		684 => "011000101100100010101",
		685 => "011000101100100010101",
		686 => "011000101100100010101",
		687 => "011000101100100010101",
		688 => "011000101100100010101",
		689 => "011000101100100010101",
		690 => "011000101100100010101",
		691 => "011000101100100010101",
		692 => "011000101100100010101",
		693 => "011000101100100010101",
		694 => "011000101100100010101",
		695 => "011000101100100010101",
		696 => "011000101100100010101",
		697 => "011000101100100010101",
		698 => "011000101100100010101",
		699 => "011000101100100010101",
		700 => "011000101100100010101",
		701 => "011000101100100010101",
		702 => "011000101100100010101",
		703 => "011000101100100010101",
		704 => "011000101100100010101",
		705 => "011000101100100010101",
		706 => "011000101100100010101",
		707 => "011000101100100010101",
		708 => "011000101100100010101",
		709 => "011000101100100010101",
		710 => "011000101100100010101",
		711 => "011000101100100010101",
		712 => "011000101100100010101",
		713 => "011000101100100010101",
		714 => "011000101100100010101",
		715 => "011000101100100010101",
		716 => "011000101100100010101",
		717 => "011000101100100010101",
		718 => "011000101100100010101",
		719 => "011000101100100010101",
		720 => "011000101100100010101",
		721 => "011000101100100010101",
		722 => "011000101100100010101",
		723 => "011000101100100010101",
		724 => "011000101100100010101",
		725 => "011000101100100010101",
		726 => "011000101100100010101",
		727 => "011000101100100010101",
		728 => "011000101100100010101",
		729 => "011000101100100010101",
		730 => "011000101100100010101",
		731 => "011000101100100010101",
		732 => "011000101100100010101",
		733 => "011000101100100010101",
		734 => "011000101100100010101",
		735 => "011000101100100010101",
		736 => "011000101100100010101",
		737 => "011000101100100010101",
		738 => "011000101100100010101",
		739 => "011000101100100010101",
		740 => "011000101100100010101",
		741 => "011000101100100010101",
		742 => "011000101100100010101",
		743 => "011000101100100010101",
		744 => "011000101100100010101",
		745 => "011000101100100010101",
		746 => "011000101100100010101",
		747 => "011000101100100010101",
		748 => "011000101100100010101",
		749 => "011000101100100010101",
		750 => "011000101100100010101",
		751 => "011000101100100010101",
		752 => "011000101100100010101",
		753 => "011000101100100010101",
		754 => "011000101100100010101",
		755 => "011000101100100010101",
		756 => "011000101100100010101",
		757 => "011000101100100010101",
		758 => "011000101100100010101",
		759 => "011000101100100010101",
		760 => "011000101100100010101",
		761 => "011000101100100010101",
		762 => "011000101100100010101",
		763 => "011000101100100010101",
		764 => "011000101100100010101",
		765 => "011000101100100010101",
		766 => "011000101100100010101",
		767 => "011000101100100010101",
		768 => "011000101100100110010",
		769 => "011000101100100110010",
		770 => "011000101100100110010",
		771 => "011000101100100110010",
		772 => "011000101100100110010",
		773 => "011000101100100110010",
		774 => "011000101100100110010",
		775 => "011000101100100110010",
		776 => "011000101100100110010",
		777 => "011000101100100110010",
		778 => "011000101100100110010",
		779 => "011000101100100110010",
		780 => "011000101100100110010",
		781 => "011000101100100110010",
		782 => "011000101100100110010",
		783 => "011000101100100110010",
		784 => "011000101100100110010",
		785 => "011000101100100110010",
		786 => "011000101100100110010",
		787 => "011000101100100110010",
		788 => "011000101100100110010",
		789 => "011000101100100110010",
		790 => "011000101100100110010",
		791 => "011000101100100110010",
		792 => "011000101100100110010",
		793 => "011000101100100110010",
		794 => "011000101100100110010",
		795 => "011000101100100110010",
		796 => "011000101100100110010",
		797 => "011000101100100110010",
		798 => "011000101100100110010",
		799 => "011000101100100110010",
		800 => "011000101100100110010",
		801 => "011000101100100110010",
		802 => "011000101100100110010",
		803 => "011000101100100110010",
		804 => "011000101100100110010",
		805 => "011000101100100110010",
		806 => "011000101100100110010",
		807 => "011000101100100110010",
		808 => "011000101100100110010",
		809 => "011000101100100110010",
		810 => "011000101100100110010",
		811 => "011000101100100110010",
		812 => "011000101100100110010",
		813 => "011000101100100110010",
		814 => "011000101100100110010",
		815 => "011000101100100110010",
		816 => "011000101100100110010",
		817 => "011000101100100110010",
		818 => "011000101100100110010",
		819 => "011000101100100110010",
		820 => "011000101100100110010",
		821 => "011000101100100110010",
		822 => "011000101100100110010",
		823 => "011000101100100110010",
		824 => "011000101100100110010",
		825 => "011000101100100110010",
		826 => "011000101100100110010",
		827 => "011000101100100110010",
		828 => "011000101100100110010",
		829 => "011000101100100110010",
		830 => "011000101100100110010",
		831 => "011000101100100110010",
		832 => "011000101100100110010",
		833 => "011000101100100110010",
		834 => "011000101100100110010",
		835 => "011000101100100110010",
		836 => "011000101100100110010",
		837 => "011000101100100110010",
		838 => "011000101100100110010",
		839 => "011000101100100110010",
		840 => "011000101100100110010",
		841 => "011000101100100110010",
		842 => "011000101100100110010",
		843 => "011000101100100110010",
		844 => "011000101100100110010",
		845 => "011000101100100110010",
		846 => "011000101100100110010",
		847 => "011000101100100110010",
		848 => "011000101100100110010",
		849 => "011000101100100110010",
		850 => "011000101100100110010",
		851 => "011000101100100110010",
		852 => "011000101100100110010",
		853 => "011000101100100110010",
		854 => "011000101100100110010",
		855 => "011000101100100110010",
		856 => "011000101100100110010",
		857 => "011000101100100110010",
		858 => "011000101100100110010",
		859 => "011000101100100110010",
		860 => "011000101100100110010",
		861 => "011000101100100110010",
		862 => "011000101100100110010",
		863 => "011000101100100110010");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;