library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT1024p_8 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT1024p_8;

architecture Behavioral of ROMFFT1024p_8 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 9 
	constant ROM_tb : ROM := (
		0 => "011000000110011110100",
		1 => "011000000110011110100",
		2 => "011000000110011110100",
		3 => "011000000101111110011",
		4 => "011000000101111110011",
		5 => "011000000101111110011",
		6 => "011000000101110011001",
		7 => "011000000101110011001",
		8 => "011000000101110011001",
		9 => "011010100100001110100",
		10 => "011010100100001110100",
		11 => "011010100100001110100",
		12 => "011000001110100010101",
		13 => "011000001110100010101",
		14 => "011000001110100010101",
		15 => "001010111100001010101",
		16 => "001010111100001010101",
		17 => "001010111100001010101",
		18 => "001001111100001010101",
		19 => "001001111100001010101",
		20 => "001001111100001010101",
		21 => "011001111100001010110",
		22 => "011001111100001010110",
		23 => "011001111100001010110",
		24 => "011000000100111010110",
		25 => "011000000100111010110",
		26 => "011000000100111010110",
		27 => "011001011101001010000",
		28 => "011001011101001010000",
		29 => "011001011101001010000",
		30 => "001011011100001010111",
		31 => "001011011100001010111",
		32 => "001011011100001010111",
		33 => "011000001101100010011",
		34 => "011000001101100010011",
		35 => "011000001101100010011",
		36 => "001001111100001010110",
		37 => "001001111100001010110",
		38 => "001001111100001010110",
		39 => "001000111100011110011",
		40 => "001000111100011110011",
		41 => "001000111100011110011",
		42 => "011001011100111010000",
		43 => "011001011100111010000",
		44 => "011001011100111010000",
		45 => "011000101100100010101",
		46 => "011000101100100010101",
		47 => "011000101100100010101",
		48 => "011001011100001010011",
		49 => "011001011100001010011",
		50 => "011001011100001010011",
		51 => "011000101100111010001",
		52 => "011000101100111010001",
		53 => "011000101100111010001",
		54 => "011000000101101010011",
		55 => "011000000101101010011",
		56 => "011000000101101010011",
		57 => "111011010100001010011",
		58 => "111011010100001010011",
		59 => "111011010100001010011",
		60 => "011000111100001010011",
		61 => "011000111100001010011",
		62 => "011000111100001010011",
		63 => "011001011100001010100",
		64 => "011001011100001010100",
		65 => "011001011100001010100",
		66 => "011000001101110010011",
		67 => "011000001101110010011",
		68 => "011000001101110010011",
		69 => "011001100100001110001",
		70 => "011001100100001110001",
		71 => "011001100100001110001",
		72 => "011000000101011010011",
		73 => "011000000101011010011",
		74 => "011000000101011010011",
		75 => "011000000101011010101",
		76 => "011000000101011010101",
		77 => "011000000101011010101",
		78 => "011000001110100010101",
		79 => "011000001110100010101",
		80 => "011000001110100010101",
		81 => "011010100100001010100",
		82 => "011010100100001010100",
		83 => "011010100100001010100",
		84 => "011000010100111010110",
		85 => "011000010100111010110",
		86 => "011000010100111010110",
		87 => "011011100100001110011",
		88 => "011011100100001110011",
		89 => "011011100100001110011",
		90 => "011000000110011010100",
		91 => "011000000110011010100",
		92 => "011000000110011010100",
		93 => "011000101100100110010",
		94 => "011000101100100110010",
		95 => "011000101100100110010",
		96 => "011000000101111110011",
		97 => "011000000101111110011",
		98 => "011000000101111110011",
		99 => "011010100100001110100",
		100 => "011010100100001110100",
		101 => "011010100100001110100",
		102 => "001010111100001010101",
		103 => "001010111100001010101",
		104 => "001010111100001010101",
		105 => "011001111100001010110",
		106 => "011001111100001010110",
		107 => "011001111100001010110",
		108 => "011001011101001010000",
		109 => "011001011101001010000",
		110 => "011001011101001010000",
		111 => "011000001101100010011",
		112 => "011000001101100010011",
		113 => "011000001101100010011",
		114 => "001000111100011110011",
		115 => "001000111100011110011",
		116 => "001000111100011110011",
		117 => "011000101100100010101",
		118 => "011000101100100010101",
		119 => "011000101100100010101",
		120 => "011000101100111010001",
		121 => "011000101100111010001",
		122 => "011000101100111010001",
		123 => "111011010100001010011",
		124 => "111011010100001010011",
		125 => "111011010100001010011",
		126 => "011001011100001010100",
		127 => "011001011100001010100",
		128 => "011001011100001010100",
		129 => "011001100100001110001",
		130 => "011001100100001110001",
		131 => "011001100100001110001",
		132 => "011000000101011010101",
		133 => "011000000101011010101",
		134 => "011000000101011010101",
		135 => "011010100100001010100",
		136 => "011010100100001010100",
		137 => "011010100100001010100",
		138 => "011011100100001110011",
		139 => "011011100100001110011",
		140 => "011011100100001110011",
		141 => "011000101100100110010",
		142 => "011000101100100110010",
		143 => "011000101100100110010",
		144 => "001001111100001010111",
		145 => "001001111100001010111",
		146 => "001001111100001010111",
		147 => "011010100100001110100",
		148 => "011010100100001110100",
		149 => "011010100100001110100",
		150 => "011010100100001010101",
		151 => "011010100100001010101",
		152 => "011010100100001010101",
		153 => "011011000100001110011",
		154 => "011011000100001110011",
		155 => "011011000100001110011",
		156 => "011010000100001010010",
		157 => "011010000100001010010",
		158 => "011010000100001010010",
		159 => "011000001101100010011",
		160 => "011000001101100010011",
		161 => "011000001101100010011",
		162 => "001000100100111010001",
		163 => "001000100100111010001",
		164 => "001000100100111010001",
		165 => "011000101100100010101",
		166 => "011000101100100010101",
		167 => "011000101100100010101",
		168 => "001000000100101110110",
		169 => "001000000100101110110",
		170 => "001000000100101110110",
		171 => "011000001101100010011",
		172 => "011000001101100010011",
		173 => "011000001101100010011",
		174 => "011010000100001110010",
		175 => "011010000100001110010",
		176 => "011010000100001110010",
		177 => "001000111100111010000",
		178 => "001000111100111010000",
		179 => "001000111100111010000",
		180 => "011000000101011010101",
		181 => "011000000101011010101",
		182 => "011000000101011010101",
		183 => "011010100100001010100",
		184 => "011010100100001010100",
		185 => "011010100100001010100",
		186 => "011000000101111010011",
		187 => "011000000101111010011",
		188 => "011000000101111010011",
		189 => "111000010100001010000",
		190 => "111000010100001010000",
		191 => "111000010100001010000",
		192 => "011010100100001110100",
		193 => "011010100100001110100",
		194 => "011010100100001110100",
		195 => "011001111100001010110",
		196 => "011001111100001010110",
		197 => "011001111100001010110",
		198 => "011000001101100010011",
		199 => "011000001101100010011",
		200 => "011000001101100010011",
		201 => "011000101100100010101",
		202 => "011000101100100010101",
		203 => "011000101100100010101",
		204 => "111011010100001010011",
		205 => "111011010100001010011",
		206 => "111011010100001010011",
		207 => "011001100100001110001",
		208 => "011001100100001110001",
		209 => "011001100100001110001",
		210 => "011010100100001010100",
		211 => "011010100100001010100",
		212 => "011010100100001010100",
		213 => "011000101100100110010",
		214 => "011000101100100110010",
		215 => "011000101100100110010",
		216 => "011010100100001110100",
		217 => "011010100100001110100",
		218 => "011010100100001110100",
		219 => "011011000100001110011",
		220 => "011011000100001110011",
		221 => "011011000100001110011",
		222 => "011000001101100010011",
		223 => "011000001101100010011",
		224 => "011000001101100010011",
		225 => "011000101100100010101",
		226 => "011000101100100010101",
		227 => "011000101100100010101",
		228 => "011000001101100010011",
		229 => "011000001101100010011",
		230 => "011000001101100010011",
		231 => "001000111100111010000",
		232 => "001000111100111010000",
		233 => "001000111100111010000",
		234 => "011010100100001010100",
		235 => "011010100100001010100",
		236 => "011010100100001010100",
		237 => "111000010100001010000",
		238 => "111000010100001010000",
		239 => "111000010100001010000",
		240 => "011010100100001110100",
		241 => "011010100100001110100",
		242 => "011010100100001110100",
		243 => "011001111100001010110",
		244 => "011001111100001010110",
		245 => "011001111100001010110",
		246 => "011000001101100010011",
		247 => "011000001101100010011",
		248 => "011000001101100010011",
		249 => "011000101100100010101",
		250 => "011000101100100010101",
		251 => "011000101100100010101",
		252 => "111011010100001010011",
		253 => "111011010100001010011",
		254 => "111011010100001010011",
		255 => "011001100100001110001",
		256 => "011001100100001110001",
		257 => "011001100100001110001",
		258 => "011010100100001010100",
		259 => "011010100100001010100",
		260 => "011010100100001010100",
		261 => "011000101100100110010",
		262 => "011000101100100110010",
		263 => "011000101100100110010",
		264 => "011010100100001110100",
		265 => "011010100100001110100",
		266 => "011010100100001110100",
		267 => "011011000100001110011",
		268 => "011011000100001110011",
		269 => "011011000100001110011",
		270 => "011000001101100010011",
		271 => "011000001101100010011",
		272 => "011000001101100010011",
		273 => "011000101100100010101",
		274 => "011000101100100010101",
		275 => "011000101100100010101",
		276 => "011000001101100010011",
		277 => "011000001101100010011",
		278 => "011000001101100010011",
		279 => "001000111100111010000",
		280 => "001000111100111010000",
		281 => "001000111100111010000",
		282 => "011010100100001010100",
		283 => "011010100100001010100",
		284 => "011010100100001010100",
		285 => "111000010100001010000",
		286 => "111000010100001010000",
		287 => "111000010100001010000",
		288 => "011001111100001010110",
		289 => "011001111100001010110",
		290 => "011001111100001010110",
		291 => "011000101100100010101",
		292 => "011000101100100010101",
		293 => "011000101100100010101",
		294 => "011001100100001110001",
		295 => "011001100100001110001",
		296 => "011001100100001110001",
		297 => "011000101100100110010",
		298 => "011000101100100110010",
		299 => "011000101100100110010",
		300 => "011011000100001110011",
		301 => "011011000100001110011",
		302 => "011011000100001110011",
		303 => "011000101100100010101",
		304 => "011000101100100010101",
		305 => "011000101100100010101",
		306 => "001000111100111010000",
		307 => "001000111100111010000",
		308 => "001000111100111010000",
		309 => "111000010100001010000",
		310 => "111000010100001010000",
		311 => "111000010100001010000",
		312 => "011001111100001010110",
		313 => "011001111100001010110",
		314 => "011001111100001010110",
		315 => "011000101100100010101",
		316 => "011000101100100010101",
		317 => "011000101100100010101",
		318 => "011001100100001110001",
		319 => "011001100100001110001",
		320 => "011001100100001110001",
		321 => "011000101100100110010",
		322 => "011000101100100110010",
		323 => "011000101100100110010",
		324 => "011011000100001110011",
		325 => "011011000100001110011",
		326 => "011011000100001110011",
		327 => "011000101100100010101",
		328 => "011000101100100010101",
		329 => "011000101100100010101",
		330 => "001000111100111010000",
		331 => "001000111100111010000",
		332 => "001000111100111010000",
		333 => "111000010100001010000",
		334 => "111000010100001010000",
		335 => "111000010100001010000",
		336 => "011001111100001010110",
		337 => "011001111100001010110",
		338 => "011001111100001010110",
		339 => "011000101100100010101",
		340 => "011000101100100010101",
		341 => "011000101100100010101",
		342 => "011001100100001110001",
		343 => "011001100100001110001",
		344 => "011001100100001110001",
		345 => "011000101100100110010",
		346 => "011000101100100110010",
		347 => "011000101100100110010",
		348 => "011011000100001110011",
		349 => "011011000100001110011",
		350 => "011011000100001110011",
		351 => "011000101100100010101",
		352 => "011000101100100010101",
		353 => "011000101100100010101",
		354 => "001000111100111010000",
		355 => "001000111100111010000",
		356 => "001000111100111010000",
		357 => "111000010100001010000",
		358 => "111000010100001010000",
		359 => "111000010100001010000",
		360 => "011001111100001010110",
		361 => "011001111100001010110",
		362 => "011001111100001010110",
		363 => "011000101100100010101",
		364 => "011000101100100010101",
		365 => "011000101100100010101",
		366 => "011001100100001110001",
		367 => "011001100100001110001",
		368 => "011001100100001110001",
		369 => "011000101100100110010",
		370 => "011000101100100110010",
		371 => "011000101100100110010",
		372 => "011011000100001110011",
		373 => "011011000100001110011",
		374 => "011011000100001110011",
		375 => "011000101100100010101",
		376 => "011000101100100010101",
		377 => "011000101100100010101",
		378 => "001000111100111010000",
		379 => "001000111100111010000",
		380 => "001000111100111010000",
		381 => "111000010100001010000",
		382 => "111000010100001010000",
		383 => "111000010100001010000",
		384 => "011000101100100010101",
		385 => "011000101100100010101",
		386 => "011000101100100010101",
		387 => "011000101100100110010",
		388 => "011000101100100110010",
		389 => "011000101100100110010",
		390 => "011000101100100010101",
		391 => "011000101100100010101",
		392 => "011000101100100010101",
		393 => "111000010100001010000",
		394 => "111000010100001010000",
		395 => "111000010100001010000",
		396 => "011000101100100010101",
		397 => "011000101100100010101",
		398 => "011000101100100010101",
		399 => "011000101100100110010",
		400 => "011000101100100110010",
		401 => "011000101100100110010",
		402 => "011000101100100010101",
		403 => "011000101100100010101",
		404 => "011000101100100010101",
		405 => "111000010100001010000",
		406 => "111000010100001010000",
		407 => "111000010100001010000",
		408 => "011000101100100010101",
		409 => "011000101100100010101",
		410 => "011000101100100010101",
		411 => "011000101100100110010",
		412 => "011000101100100110010",
		413 => "011000101100100110010",
		414 => "011000101100100010101",
		415 => "011000101100100010101",
		416 => "011000101100100010101",
		417 => "111000010100001010000",
		418 => "111000010100001010000",
		419 => "111000010100001010000",
		420 => "011000101100100010101",
		421 => "011000101100100010101",
		422 => "011000101100100010101",
		423 => "011000101100100110010",
		424 => "011000101100100110010",
		425 => "011000101100100110010",
		426 => "011000101100100010101",
		427 => "011000101100100010101",
		428 => "011000101100100010101",
		429 => "111000010100001010000",
		430 => "111000010100001010000",
		431 => "111000010100001010000",
		432 => "011000101100100010101",
		433 => "011000101100100010101",
		434 => "011000101100100010101",
		435 => "011000101100100110010",
		436 => "011000101100100110010",
		437 => "011000101100100110010",
		438 => "011000101100100010101",
		439 => "011000101100100010101",
		440 => "011000101100100010101",
		441 => "111000010100001010000",
		442 => "111000010100001010000",
		443 => "111000010100001010000",
		444 => "011000101100100010101",
		445 => "011000101100100010101",
		446 => "011000101100100010101",
		447 => "011000101100100110010",
		448 => "011000101100100110010",
		449 => "011000101100100110010",
		450 => "011000101100100010101",
		451 => "011000101100100010101",
		452 => "011000101100100010101",
		453 => "111000010100001010000",
		454 => "111000010100001010000",
		455 => "111000010100001010000",
		456 => "011000101100100010101",
		457 => "011000101100100010101",
		458 => "011000101100100010101",
		459 => "011000101100100110010",
		460 => "011000101100100110010",
		461 => "011000101100100110010",
		462 => "011000101100100010101",
		463 => "011000101100100010101",
		464 => "011000101100100010101",
		465 => "111000010100001010000",
		466 => "111000010100001010000",
		467 => "111000010100001010000",
		468 => "011000101100100010101",
		469 => "011000101100100010101",
		470 => "011000101100100010101",
		471 => "011000101100100110010",
		472 => "011000101100100110010",
		473 => "011000101100100110010",
		474 => "011000101100100010101",
		475 => "011000101100100010101",
		476 => "011000101100100010101",
		477 => "111000010100001010000",
		478 => "111000010100001010000",
		479 => "111000010100001010000",
		480 => "011000101100100110010",
		481 => "011000101100100110010",
		482 => "011000101100100110010",
		483 => "111000010100001010000",
		484 => "111000010100001010000",
		485 => "111000010100001010000",
		486 => "011000101100100110010",
		487 => "011000101100100110010",
		488 => "011000101100100110010",
		489 => "111000010100001010000",
		490 => "111000010100001010000",
		491 => "111000010100001010000",
		492 => "011000101100100110010",
		493 => "011000101100100110010",
		494 => "011000101100100110010",
		495 => "111000010100001010000",
		496 => "111000010100001010000",
		497 => "111000010100001010000",
		498 => "011000101100100110010",
		499 => "011000101100100110010",
		500 => "011000101100100110010",
		501 => "111000010100001010000",
		502 => "111000010100001010000",
		503 => "111000010100001010000",
		504 => "011000101100100110010",
		505 => "011000101100100110010",
		506 => "011000101100100110010",
		507 => "111000010100001010000",
		508 => "111000010100001010000",
		509 => "111000010100001010000",
		510 => "011000101100100110010",
		511 => "011000101100100110010",
		512 => "011000101100100110010",
		513 => "111000010100001010000",
		514 => "111000010100001010000",
		515 => "111000010100001010000",
		516 => "011000101100100110010",
		517 => "011000101100100110010",
		518 => "011000101100100110010",
		519 => "111000010100001010000",
		520 => "111000010100001010000",
		521 => "111000010100001010000",
		522 => "011000101100100110010",
		523 => "011000101100100110010",
		524 => "011000101100100110010",
		525 => "111000010100001010000",
		526 => "111000010100001010000",
		527 => "111000010100001010000",
		528 => "011000101100100110010",
		529 => "011000101100100110010",
		530 => "011000101100100110010",
		531 => "111000010100001010000",
		532 => "111000010100001010000",
		533 => "111000010100001010000",
		534 => "011000101100100110010",
		535 => "011000101100100110010",
		536 => "011000101100100110010",
		537 => "111000010100001010000",
		538 => "111000010100001010000",
		539 => "111000010100001010000",
		540 => "011000101100100110010",
		541 => "011000101100100110010",
		542 => "011000101100100110010",
		543 => "111000010100001010000",
		544 => "111000010100001010000",
		545 => "111000010100001010000",
		546 => "011000101100100110010",
		547 => "011000101100100110010",
		548 => "011000101100100110010",
		549 => "111000010100001010000",
		550 => "111000010100001010000",
		551 => "111000010100001010000",
		552 => "011000101100100110010",
		553 => "011000101100100110010",
		554 => "011000101100100110010",
		555 => "111000010100001010000",
		556 => "111000010100001010000",
		557 => "111000010100001010000",
		558 => "011000101100100110010",
		559 => "011000101100100110010",
		560 => "011000101100100110010",
		561 => "111000010100001010000",
		562 => "111000010100001010000",
		563 => "111000010100001010000",
		564 => "011000101100100110010",
		565 => "011000101100100110010",
		566 => "011000101100100110010",
		567 => "111000010100001010000",
		568 => "111000010100001010000",
		569 => "111000010100001010000",
		570 => "011000101100100110010",
		571 => "011000101100100110010",
		572 => "011000101100100110010",
		573 => "111000010100001010000",
		574 => "111000010100001010000",
		575 => "111000010100001010000",
		576 => "111000010100001010000",
		577 => "111000010100001010000",
		578 => "111000010100001010000",
		579 => "111000010100001010000",
		580 => "111000010100001010000",
		581 => "111000010100001010000",
		582 => "111000010100001010000",
		583 => "111000010100001010000",
		584 => "111000010100001010000",
		585 => "111000010100001010000",
		586 => "111000010100001010000",
		587 => "111000010100001010000",
		588 => "111000010100001010000",
		589 => "111000010100001010000",
		590 => "111000010100001010000",
		591 => "111000010100001010000",
		592 => "111000010100001010000",
		593 => "111000010100001010000",
		594 => "111000010100001010000",
		595 => "111000010100001010000",
		596 => "111000010100001010000",
		597 => "111000010100001010000",
		598 => "111000010100001010000",
		599 => "111000010100001010000",
		600 => "111000010100001010000",
		601 => "111000010100001010000",
		602 => "111000010100001010000",
		603 => "111000010100001010000",
		604 => "111000010100001010000",
		605 => "111000010100001010000",
		606 => "111000010100001010000",
		607 => "111000010100001010000",
		608 => "111000010100001010000",
		609 => "111000010100001010000",
		610 => "111000010100001010000",
		611 => "111000010100001010000",
		612 => "111000010100001010000",
		613 => "111000010100001010000",
		614 => "111000010100001010000",
		615 => "111000010100001010000",
		616 => "111000010100001010000",
		617 => "111000010100001010000",
		618 => "111000010100001010000",
		619 => "111000010100001010000",
		620 => "111000010100001010000",
		621 => "111000010100001010000",
		622 => "111000010100001010000",
		623 => "111000010100001010000",
		624 => "111000010100001010000",
		625 => "111000010100001010000",
		626 => "111000010100001010000",
		627 => "111000010100001010000",
		628 => "111000010100001010000",
		629 => "111000010100001010000",
		630 => "111000010100001010000",
		631 => "111000010100001010000",
		632 => "111000010100001010000",
		633 => "111000010100001010000",
		634 => "111000010100001010000",
		635 => "111000010100001010000",
		636 => "111000010100001010000",
		637 => "111000010100001010000",
		638 => "111000010100001010000",
		639 => "111000010100001010000",
		640 => "111000010100001010000",
		641 => "111000010100001010000",
		642 => "111000010100001010000",
		643 => "111000010100001010000",
		644 => "111000010100001010000",
		645 => "111000010100001010000",
		646 => "111000010100001010000",
		647 => "111000010100001010000",
		648 => "111000010100001010000",
		649 => "111000010100001010000",
		650 => "111000010100001010000",
		651 => "111000010100001010000",
		652 => "111000010100001010000",
		653 => "111000010100001010000",
		654 => "111000010100001010000",
		655 => "111000010100001010000",
		656 => "111000010100001010000",
		657 => "111000010100001010000",
		658 => "111000010100001010000",
		659 => "111000010100001010000",
		660 => "111000010100001010000",
		661 => "111000010100001010000",
		662 => "111000010100001010000",
		663 => "111000010100001010000",
		664 => "111000010100001010000",
		665 => "111000010100001010000",
		666 => "111000010100001010000",
		667 => "111000010100001010000",
		668 => "111000010100001010000",
		669 => "111000010100001010000",
		670 => "111000010100001010000",
		671 => "111000010100001010000",
		672 => "111000010100001010000",
		673 => "111000010100001010000",
		674 => "111000010100001010000",
		675 => "111000010100001010000",
		676 => "111000010100001010000",
		677 => "111000010100001010000",
		678 => "111000010100001010000",
		679 => "111000010100001010000",
		680 => "111000010100001010000",
		681 => "111000010100001010000",
		682 => "111000010100001010000",
		683 => "111000010100001010000",
		684 => "111000010100001010000",
		685 => "111000010100001010000",
		686 => "111000010100001010000",
		687 => "111000010100001010000",
		688 => "111000010100001010000",
		689 => "111000010100001010000",
		690 => "111000010100001010000",
		691 => "111000010100001010000",
		692 => "111000010100001010000",
		693 => "111000010100001010000",
		694 => "111000010100001010000",
		695 => "111000010100001010000",
		696 => "111000010100001010000",
		697 => "111000010100001010000",
		698 => "111000010100001010000",
		699 => "111000010100001010000",
		700 => "111000010100001010000",
		701 => "111000010100001010000",
		702 => "111000010100001010000",
		703 => "111000010100001010000",
		704 => "111000010100001010000",
		705 => "111000010100001010000",
		706 => "111000010100001010000",
		707 => "111000010100001010000",
		708 => "111000010100001010000",
		709 => "111000010100001010000",
		710 => "111000010100001010000",
		711 => "111000010100001010000",
		712 => "111000010100001010000",
		713 => "111000010100001010000",
		714 => "111000010100001010000",
		715 => "111000010100001010000",
		716 => "111000010100001010000",
		717 => "111000010100001010000",
		718 => "111000010100001010000",
		719 => "111000010100001010000",
		720 => "111000010100001010000",
		721 => "111000010100001010000",
		722 => "111000010100001010000",
		723 => "111000010100001010000",
		724 => "111000010100001010000",
		725 => "111000010100001010000",
		726 => "111000010100001010000",
		727 => "111000010100001010000",
		728 => "111000010100001010000",
		729 => "111000010100001010000",
		730 => "111000010100001010000",
		731 => "111000010100001010000",
		732 => "111000010100001010000",
		733 => "111000010100001010000",
		734 => "111000010100001010000",
		735 => "111000010100001010000",
		736 => "111000010100001010000",
		737 => "111000010100001010000",
		738 => "111000010100001010000",
		739 => "111000010100001010000",
		740 => "111000010100001010000",
		741 => "111000010100001010000",
		742 => "111000010100001010000",
		743 => "111000010100001010000",
		744 => "111000010100001010000",
		745 => "111000010100001010000",
		746 => "111000010100001010000",
		747 => "111000010100001010000",
		748 => "111000010100001010000",
		749 => "111000010100001010000",
		750 => "111000010100001010000",
		751 => "111000010100001010000",
		752 => "111000010100001010000",
		753 => "111000010100001010000",
		754 => "111000010100001010000",
		755 => "111000010100001010000",
		756 => "111000010100001010000",
		757 => "111000010100001010000",
		758 => "111000010100001010000",
		759 => "111000010100001010000",
		760 => "111000010100001010000",
		761 => "111000010100001010000",
		762 => "111000010100001010000",
		763 => "111000010100001010000",
		764 => "111000010100001010000",
		765 => "111000010100001010000",
		766 => "111000010100001010000",
		767 => "111000010100001010000",
		768 => "111000010100001010000",
		769 => "111000010100001010000",
		770 => "111000010100001010000",
		771 => "111000010100001010000",
		772 => "111000010100001010000",
		773 => "111000010100001010000",
		774 => "111000010100001010000",
		775 => "111000010100001010000",
		776 => "111000010100001010000",
		777 => "111000010100001010000",
		778 => "111000010100001010000",
		779 => "111000010100001010000",
		780 => "111000010100001010000",
		781 => "111000010100001010000",
		782 => "111000010100001010000",
		783 => "111000010100001010000",
		784 => "111000010100001010000",
		785 => "111000010100001010000",
		786 => "111000010100001010000",
		787 => "111000010100001010000",
		788 => "111000010100001010000",
		789 => "111000010100001010000",
		790 => "111000010100001010000",
		791 => "111000010100001010000",
		792 => "111000010100001010000",
		793 => "111000010100001010000",
		794 => "111000010100001010000",
		795 => "111000010100001010000",
		796 => "111000010100001010000",
		797 => "111000010100001010000",
		798 => "111000010100001010000",
		799 => "111000010100001010000",
		800 => "111000010100001010000",
		801 => "111000010100001010000",
		802 => "111000010100001010000",
		803 => "111000010100001010000",
		804 => "111000010100001010000",
		805 => "111000010100001010000",
		806 => "111000010100001010000",
		807 => "111000010100001010000",
		808 => "111000010100001010000",
		809 => "111000010100001010000",
		810 => "111000010100001010000",
		811 => "111000010100001010000",
		812 => "111000010100001010000",
		813 => "111000010100001010000",
		814 => "111000010100001010000",
		815 => "111000010100001010000",
		816 => "111000010100001010000",
		817 => "111000010100001010000",
		818 => "111000010100001010000",
		819 => "111000010100001010000",
		820 => "111000010100001010000",
		821 => "111000010100001010000",
		822 => "111000010100001010000",
		823 => "111000010100001010000",
		824 => "111000010100001010000",
		825 => "111000010100001010000",
		826 => "111000010100001010000",
		827 => "111000010100001010000",
		828 => "111000010100001010000",
		829 => "111000010100001010000",
		830 => "111000010100001010000",
		831 => "111000010100001010000",
		832 => "111000010100001010000",
		833 => "111000010100001010000",
		834 => "111000010100001010000",
		835 => "111000010100001010000",
		836 => "111000010100001010000",
		837 => "111000010100001010000",
		838 => "111000010100001010000",
		839 => "111000010100001010000",
		840 => "111000010100001010000",
		841 => "111000010100001010000",
		842 => "111000010100001010000",
		843 => "111000010100001010000",
		844 => "111000010100001010000",
		845 => "111000010100001010000",
		846 => "111000010100001010000",
		847 => "111000010100001010000",
		848 => "111000010100001010000",
		849 => "111000010100001010000",
		850 => "111000010100001010000",
		851 => "111000010100001010000",
		852 => "111000010100001010000",
		853 => "111000010100001010000",
		854 => "111000010100001010000",
		855 => "111000010100001010000",
		856 => "111000010100001010000",
		857 => "111000010100001010000",
		858 => "111000010100001010000",
		859 => "111000010100001010000",
		860 => "111000010100001010000",
		861 => "111000010100001010000",
		862 => "111000010100001010000",
		863 => "111000010100001010000");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;