library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT3 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT3;

architecture Behavioral of ROMFFT3 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 4 
	constant ROM_tb : ROM := (
		0 => "001000011110101011000",
		1 => "001000011110101011000",
		2 => "001000011110101011000",
		3 => "011011100100001110111",
		4 => "011011100100001110111",
		5 => "011011100100001110111",
		6 => "001000000100111010010",
		7 => "001000000100111010010",
		8 => "001000000100111010010",
		9 => "011010011101011010000",
		10 => "011010011101011010000",
		11 => "011010011101011010000",
		12 => "011000000100111110001",
		13 => "011000000100111110001",
		14 => "011000000100111110001",
		15 => "011010000100001010010",
		16 => "011010000100001010010",
		17 => "011010000100001010010",
		18 => "011001001100111010000",
		19 => "011001001100111010000",
		20 => "011001001100111010000",
		21 => "011000110100011010011",
		22 => "011000110100011010011",
		23 => "011000110100011010011",
		24 => "011001100100001110000",
		25 => "011001100100001110000",
		26 => "011001100100001110000",
		27 => "001000100100111110001",
		28 => "001000100100111110001",
		29 => "001000100100111110001",
		30 => "011001000100001110001",
		31 => "011001000100001110001",
		32 => "011001000100001110001",
		33 => "011001011100001010100",
		34 => "011001011100001010100",
		35 => "011001011100001010100",
		36 => "011000000101111010010",
		37 => "011000000101111010010",
		38 => "011000000101111010010",
		39 => "011000000101011010101",
		40 => "011000000101011010101",
		41 => "011000000101011010101",
		42 => "011000000101111010011",
		43 => "011000000101111010011",
		44 => "011000000101111010011",
		45 => "011000000110011010110",
		46 => "011000000110011010110",
		47 => "011000000110011010110",
		48 => "001000011110101011000",
		49 => "001000011110101011000",
		50 => "001000011110101011000",
		51 => "011000001111010010111",
		52 => "011000001111010010111",
		53 => "011000001111010010111",
		54 => "001000000100111010010",
		55 => "001000000100111010010",
		56 => "001000000100111010010",
		57 => "011010100100001010100",
		58 => "011010100100001010100",
		59 => "011010100100001010100",
		60 => "001000111100001010011",
		61 => "001000111100001010011",
		62 => "001000111100001010011",
		63 => "011001011101001010000",
		64 => "011001011101001010000",
		65 => "011001011101001010000",
		66 => "001000011100111010001",
		67 => "001000011100111010001",
		68 => "001000011100111010001",
		69 => "011000110100011010011",
		70 => "011000110100011010011",
		71 => "011000110100011010011",
		72 => "001000011100111010000",
		73 => "001000011100111010000",
		74 => "001000011100111010000",
		75 => "001000110100011010011",
		76 => "001000110100011010011",
		77 => "001000110100011010011",
		78 => "011001000100001110001",
		79 => "011001000100001110001",
		80 => "011001000100001110001",
		81 => "011010000100001110010",
		82 => "011010000100001110010",
		83 => "011010000100001110010",
		84 => "011000000101111010010",
		85 => "011000000101111010010",
		86 => "011000000101111010010",
		87 => "011000001110100010101",
		88 => "011000001110100010101",
		89 => "011000001110100010101",
		90 => "001001111101111010000",
		91 => "001001111101111010000",
		92 => "001001111101111010000",
		93 => "001000011101001111001",
		94 => "001000011101001111001",
		95 => "001000011101001111001",
		96 => "011100001110011010000",
		97 => "011100001110011010000",
		98 => "011100001110011010000",
		99 => "001001011100001010110",
		100 => "001001011100001010110",
		101 => "001001011100001010110",
		102 => "001000011100111010001",
		103 => "001000011100111010001",
		104 => "001000011100111010001",
		105 => "011000000100111010000",
		106 => "011000000100111010000",
		107 => "011000000100111010000",
		108 => "011000000100111010010",
		109 => "011000000100111010010",
		110 => "011000000100111010010",
		111 => "011000000101001010001",
		112 => "011000000101001010001",
		113 => "011000000101001010001",
		114 => "001000011100101110011",
		115 => "001000011100101110011",
		116 => "001000011100101110011",
		117 => "011000000101111010011",
		118 => "011000000101111010011",
		119 => "011000000101111010011",
		120 => "001000011110011010111",
		121 => "001000011110011010111",
		122 => "001000011110011010111",
		123 => "011011000100001010010",
		124 => "011011000100001010010",
		125 => "011011000100001010010",
		126 => "011010000100001010100",
		127 => "011010000100001010100",
		128 => "011010000100001010100",
		129 => "011001100100001110000",
		130 => "011001100100001110000",
		131 => "011001100100001110000",
		132 => "011000000101101010001",
		133 => "011000000101101010001",
		134 => "011000000101101010001",
		135 => "011000000101001010001",
		136 => "011000000101001010001",
		137 => "011000000101001010001",
		138 => "011001100100011010000",
		139 => "011001100100011010000",
		140 => "011001100100011010000",
		141 => "001001111101111010000",
		142 => "001001111101111010000",
		143 => "001001111101111010000",
		144 => "011100001110011010000",
		145 => "011100001110011010000",
		146 => "011100001110011010000",
		147 => "001001011100001010110",
		148 => "001001011100001010110",
		149 => "001001011100001010110",
		150 => "001000011100111010001",
		151 => "001000011100111010001",
		152 => "001000011100111010001",
		153 => "011000000100111010000",
		154 => "011000000100111010000",
		155 => "011000000100111010000",
		156 => "011000000100111010010",
		157 => "011000000100111010010",
		158 => "011000000100111010010",
		159 => "011000000101001010001",
		160 => "011000000101001010001",
		161 => "011000000101001010001",
		162 => "001000011100101110011",
		163 => "001000011100101110011",
		164 => "001000011100101110011",
		165 => "011000000101111010011",
		166 => "011000000101111010011",
		167 => "011000000101111010011",
		168 => "001000011110011010111",
		169 => "001000011110011010111",
		170 => "001000011110011010111",
		171 => "011011000100001010010",
		172 => "011011000100001010010",
		173 => "011011000100001010010",
		174 => "011010000100001010100",
		175 => "011010000100001010100",
		176 => "011010000100001010100",
		177 => "011001100100001110000",
		178 => "011001100100001110000",
		179 => "011001100100001110000",
		180 => "011000000101101010001",
		181 => "011000000101101010001",
		182 => "011000000101101010001",
		183 => "011000000101001010001",
		184 => "011000000101001010001",
		185 => "011000000101001010001",
		186 => "011001100100011010000",
		187 => "011001100100011010000",
		188 => "011001100100011010000",
		189 => "001001111101111010000",
		190 => "001001111101111010000",
		191 => "001001111101111010000",
		192 => "011011101110001010000",
		193 => "011011101110001010000",
		194 => "011011101110001010000",
		195 => "011000001101100010011",
		196 => "011000001101100010011",
		197 => "011000001101100010011",
		198 => "011000101100101010100",
		199 => "011000101100101010100",
		200 => "011000101100101010100",
		201 => "011000000101011010010",
		202 => "011000000101011010010",
		203 => "011000000101011010010",
		204 => "001000011110001010110",
		205 => "001000011110001010110",
		206 => "001000011110001010110",
		207 => "011000001101100010011",
		208 => "011000001101100010011",
		209 => "011000001101100010011",
		210 => "011001000100001110100",
		211 => "011001000100001110100",
		212 => "011001000100001110100",
		213 => "011000000101011010010",
		214 => "011000000101011010010",
		215 => "011000000101011010010",
		216 => "011011101110001010000",
		217 => "011011101110001010000",
		218 => "011011101110001010000",
		219 => "011000001101100010011",
		220 => "011000001101100010011",
		221 => "011000001101100010011",
		222 => "011000101100101010100",
		223 => "011000101100101010100",
		224 => "011000101100101010100",
		225 => "011000000101011010010",
		226 => "011000000101011010010",
		227 => "011000000101011010010",
		228 => "001000011110001010110",
		229 => "001000011110001010110",
		230 => "001000011110001010110",
		231 => "011000001101100010011",
		232 => "011000001101100010011",
		233 => "011000001101100010011",
		234 => "011001000100001110100",
		235 => "011001000100001110100",
		236 => "011001000100001110100",
		237 => "011000000101011010010",
		238 => "011000000101011010010",
		239 => "011000000101011010010",
		240 => "011011101110001010000",
		241 => "011011101110001010000",
		242 => "011011101110001010000",
		243 => "011000001101100010011",
		244 => "011000001101100010011",
		245 => "011000001101100010011",
		246 => "011000101100101010100",
		247 => "011000101100101010100",
		248 => "011000101100101010100",
		249 => "011000000101011010010",
		250 => "011000000101011010010",
		251 => "011000000101011010010",
		252 => "001000011110001010110",
		253 => "001000011110001010110",
		254 => "001000011110001010110",
		255 => "011000001101100010011",
		256 => "011000001101100010011",
		257 => "011000001101100010011",
		258 => "011001000100001110100",
		259 => "011001000100001110100",
		260 => "011001000100001110100",
		261 => "011000000101011010010",
		262 => "011000000101011010010",
		263 => "011000000101011010010",
		264 => "011011101110001010000",
		265 => "011011101110001010000",
		266 => "011011101110001010000",
		267 => "011000001101100010011",
		268 => "011000001101100010011",
		269 => "011000001101100010011",
		270 => "011000101100101010100",
		271 => "011000101100101010100",
		272 => "011000101100101010100",
		273 => "011000000101011010010",
		274 => "011000000101011010010",
		275 => "011000000101011010010",
		276 => "001000011110001010110",
		277 => "001000011110001010110",
		278 => "001000011110001010110",
		279 => "011000001101100010011",
		280 => "011000001101100010011",
		281 => "011000001101100010011",
		282 => "011001000100001110100",
		283 => "011001000100001110100",
		284 => "011001000100001110100",
		285 => "011000000101011010010",
		286 => "011000000101011010010",
		287 => "011000000101011010010",
		288 => "011000000101110011001",
		289 => "011000000101110011001",
		290 => "011000000101110011001",
		291 => "011000000101101010011",
		292 => "011000000101101010011",
		293 => "011000000101101010011",
		294 => "011000000101110011001",
		295 => "011000000101110011001",
		296 => "011000000101110011001",
		297 => "011000000101101010011",
		298 => "011000000101101010011",
		299 => "011000000101101010011",
		300 => "011000000101110011001",
		301 => "011000000101110011001",
		302 => "011000000101110011001",
		303 => "011000000101101010011",
		304 => "011000000101101010011",
		305 => "011000000101101010011",
		306 => "011000000101110011001",
		307 => "011000000101110011001",
		308 => "011000000101110011001",
		309 => "011000000101101010011",
		310 => "011000000101101010011",
		311 => "011000000101101010011",
		312 => "011000000101110011001",
		313 => "011000000101110011001",
		314 => "011000000101110011001",
		315 => "011000000101101010011",
		316 => "011000000101101010011",
		317 => "011000000101101010011",
		318 => "011000000101110011001",
		319 => "011000000101110011001",
		320 => "011000000101110011001",
		321 => "011000000101101010011",
		322 => "011000000101101010011",
		323 => "011000000101101010011",
		324 => "011000000101110011001",
		325 => "011000000101110011001",
		326 => "011000000101110011001",
		327 => "011000000101101010011",
		328 => "011000000101101010011",
		329 => "011000000101101010011",
		330 => "011000000101110011001",
		331 => "011000000101110011001",
		332 => "011000000101110011001",
		333 => "011000000101101010011",
		334 => "011000000101101010011",
		335 => "011000000101101010011",
		336 => "011000000101110011001",
		337 => "011000000101110011001",
		338 => "011000000101110011001",
		339 => "011000000101101010011",
		340 => "011000000101101010011",
		341 => "011000000101101010011",
		342 => "011000000101110011001",
		343 => "011000000101110011001",
		344 => "011000000101110011001",
		345 => "011000000101101010011",
		346 => "011000000101101010011",
		347 => "011000000101101010011",
		348 => "011000000101110011001",
		349 => "011000000101110011001",
		350 => "011000000101110011001",
		351 => "011000000101101010011",
		352 => "011000000101101010011",
		353 => "011000000101101010011",
		354 => "011000000101110011001",
		355 => "011000000101110011001",
		356 => "011000000101110011001",
		357 => "011000000101101010011",
		358 => "011000000101101010011",
		359 => "011000000101101010011",
		360 => "011000000101110011001",
		361 => "011000000101110011001",
		362 => "011000000101110011001",
		363 => "011000000101101010011",
		364 => "011000000101101010011",
		365 => "011000000101101010011",
		366 => "011000000101110011001",
		367 => "011000000101110011001",
		368 => "011000000101110011001",
		369 => "011000000101101010011",
		370 => "011000000101101010011",
		371 => "011000000101101010011",
		372 => "011000000101110011001",
		373 => "011000000101110011001",
		374 => "011000000101110011001",
		375 => "011000000101101010011",
		376 => "011000000101101010011",
		377 => "011000000101101010011",
		378 => "011000000101110011001",
		379 => "011000000101110011001",
		380 => "011000000101110011001",
		381 => "011000000101101010011",
		382 => "011000000101101010011",
		383 => "011000000101101010011",
		384 => "001010111100001010101",
		385 => "001010111100001010101",
		386 => "001010111100001010101",
		387 => "011010100100001010101",
		388 => "011010100100001010101",
		389 => "011010100100001010101",
		390 => "001010111100001010101",
		391 => "001010111100001010101",
		392 => "001010111100001010101",
		393 => "011010100100001010101",
		394 => "011010100100001010101",
		395 => "011010100100001010101",
		396 => "001010111100001010101",
		397 => "001010111100001010101",
		398 => "001010111100001010101",
		399 => "011010100100001010101",
		400 => "011010100100001010101",
		401 => "011010100100001010101",
		402 => "001010111100001010101",
		403 => "001010111100001010101",
		404 => "001010111100001010101",
		405 => "011010100100001010101",
		406 => "011010100100001010101",
		407 => "011010100100001010101",
		408 => "001010111100001010101",
		409 => "001010111100001010101",
		410 => "001010111100001010101",
		411 => "011010100100001010101",
		412 => "011010100100001010101",
		413 => "011010100100001010101",
		414 => "001010111100001010101",
		415 => "001010111100001010101",
		416 => "001010111100001010101",
		417 => "011010100100001010101",
		418 => "011010100100001010101",
		419 => "011010100100001010101",
		420 => "001010111100001010101",
		421 => "001010111100001010101",
		422 => "001010111100001010101",
		423 => "011010100100001010101",
		424 => "011010100100001010101",
		425 => "011010100100001010101",
		426 => "001010111100001010101",
		427 => "001010111100001010101",
		428 => "001010111100001010101",
		429 => "011010100100001010101",
		430 => "011010100100001010101",
		431 => "011010100100001010101",
		432 => "001010111100001010101",
		433 => "001010111100001010101",
		434 => "001010111100001010101",
		435 => "011010100100001010101",
		436 => "011010100100001010101",
		437 => "011010100100001010101",
		438 => "001010111100001010101",
		439 => "001010111100001010101",
		440 => "001010111100001010101",
		441 => "011010100100001010101",
		442 => "011010100100001010101",
		443 => "011010100100001010101",
		444 => "001010111100001010101",
		445 => "001010111100001010101",
		446 => "001010111100001010101",
		447 => "011010100100001010101",
		448 => "011010100100001010101",
		449 => "011010100100001010101",
		450 => "001010111100001010101",
		451 => "001010111100001010101",
		452 => "001010111100001010101",
		453 => "011010100100001010101",
		454 => "011010100100001010101",
		455 => "011010100100001010101",
		456 => "001010111100001010101",
		457 => "001010111100001010101",
		458 => "001010111100001010101",
		459 => "011010100100001010101",
		460 => "011010100100001010101",
		461 => "011010100100001010101",
		462 => "001010111100001010101",
		463 => "001010111100001010101",
		464 => "001010111100001010101",
		465 => "011010100100001010101",
		466 => "011010100100001010101",
		467 => "011010100100001010101",
		468 => "001010111100001010101",
		469 => "001010111100001010101",
		470 => "001010111100001010101",
		471 => "011010100100001010101",
		472 => "011010100100001010101",
		473 => "011010100100001010101",
		474 => "001010111100001010101",
		475 => "001010111100001010101",
		476 => "001010111100001010101",
		477 => "011010100100001010101",
		478 => "011010100100001010101",
		479 => "011010100100001010101",
		480 => "011000001101100010011",
		481 => "011000001101100010011",
		482 => "011000001101100010011",
		483 => "011000001101100010011",
		484 => "011000001101100010011",
		485 => "011000001101100010011",
		486 => "011000001101100010011",
		487 => "011000001101100010011",
		488 => "011000001101100010011",
		489 => "011000001101100010011",
		490 => "011000001101100010011",
		491 => "011000001101100010011",
		492 => "011000001101100010011",
		493 => "011000001101100010011",
		494 => "011000001101100010011",
		495 => "011000001101100010011",
		496 => "011000001101100010011",
		497 => "011000001101100010011",
		498 => "011000001101100010011",
		499 => "011000001101100010011",
		500 => "011000001101100010011",
		501 => "011000001101100010011",
		502 => "011000001101100010011",
		503 => "011000001101100010011",
		504 => "011000001101100010011",
		505 => "011000001101100010011",
		506 => "011000001101100010011",
		507 => "011000001101100010011",
		508 => "011000001101100010011",
		509 => "011000001101100010011",
		510 => "011000001101100010011",
		511 => "011000001101100010011",
		512 => "011000001101100010011",
		513 => "011000001101100010011",
		514 => "011000001101100010011",
		515 => "011000001101100010011",
		516 => "011000001101100010011",
		517 => "011000001101100010011",
		518 => "011000001101100010011",
		519 => "011000001101100010011",
		520 => "011000001101100010011",
		521 => "011000001101100010011",
		522 => "011000001101100010011",
		523 => "011000001101100010011",
		524 => "011000001101100010011",
		525 => "011000001101100010011",
		526 => "011000001101100010011",
		527 => "011000001101100010011",
		528 => "011000001101100010011",
		529 => "011000001101100010011",
		530 => "011000001101100010011",
		531 => "011000001101100010011",
		532 => "011000001101100010011",
		533 => "011000001101100010011",
		534 => "011000001101100010011",
		535 => "011000001101100010011",
		536 => "011000001101100010011",
		537 => "011000001101100010011",
		538 => "011000001101100010011",
		539 => "011000001101100010011",
		540 => "011000001101100010011",
		541 => "011000001101100010011",
		542 => "011000001101100010011",
		543 => "011000001101100010011",
		544 => "011000001101100010011",
		545 => "011000001101100010011",
		546 => "011000001101100010011",
		547 => "011000001101100010011",
		548 => "011000001101100010011",
		549 => "011000001101100010011",
		550 => "011000001101100010011",
		551 => "011000001101100010011",
		552 => "011000001101100010011",
		553 => "011000001101100010011",
		554 => "011000001101100010011",
		555 => "011000001101100010011",
		556 => "011000001101100010011",
		557 => "011000001101100010011",
		558 => "011000001101100010011",
		559 => "011000001101100010011",
		560 => "011000001101100010011",
		561 => "011000001101100010011",
		562 => "011000001101100010011",
		563 => "011000001101100010011",
		564 => "011000001101100010011",
		565 => "011000001101100010011",
		566 => "011000001101100010011",
		567 => "011000001101100010011",
		568 => "011000001101100010011",
		569 => "011000001101100010011",
		570 => "011000001101100010011",
		571 => "011000001101100010011",
		572 => "011000001101100010011",
		573 => "011000001101100010011",
		574 => "011000001101100010011",
		575 => "011000001101100010011",
		576 => "011001100100001110001",
		577 => "011001100100001110001",
		578 => "011001100100001110001",
		579 => "011001100100001110001",
		580 => "011001100100001110001",
		581 => "011001100100001110001",
		582 => "011001100100001110001",
		583 => "011001100100001110001",
		584 => "011001100100001110001",
		585 => "011001100100001110001",
		586 => "011001100100001110001",
		587 => "011001100100001110001",
		588 => "011001100100001110001",
		589 => "011001100100001110001",
		590 => "011001100100001110001",
		591 => "011001100100001110001",
		592 => "011001100100001110001",
		593 => "011001100100001110001",
		594 => "011001100100001110001",
		595 => "011001100100001110001",
		596 => "011001100100001110001",
		597 => "011001100100001110001",
		598 => "011001100100001110001",
		599 => "011001100100001110001",
		600 => "011001100100001110001",
		601 => "011001100100001110001",
		602 => "011001100100001110001",
		603 => "011001100100001110001",
		604 => "011001100100001110001",
		605 => "011001100100001110001",
		606 => "011001100100001110001",
		607 => "011001100100001110001",
		608 => "011001100100001110001",
		609 => "011001100100001110001",
		610 => "011001100100001110001",
		611 => "011001100100001110001",
		612 => "011001100100001110001",
		613 => "011001100100001110001",
		614 => "011001100100001110001",
		615 => "011001100100001110001",
		616 => "011001100100001110001",
		617 => "011001100100001110001",
		618 => "011001100100001110001",
		619 => "011001100100001110001",
		620 => "011001100100001110001",
		621 => "011001100100001110001",
		622 => "011001100100001110001",
		623 => "011001100100001110001",
		624 => "011001100100001110001",
		625 => "011001100100001110001",
		626 => "011001100100001110001",
		627 => "011001100100001110001",
		628 => "011001100100001110001",
		629 => "011001100100001110001",
		630 => "011001100100001110001",
		631 => "011001100100001110001",
		632 => "011001100100001110001",
		633 => "011001100100001110001",
		634 => "011001100100001110001",
		635 => "011001100100001110001",
		636 => "011001100100001110001",
		637 => "011001100100001110001",
		638 => "011001100100001110001",
		639 => "011001100100001110001",
		640 => "011001100100001110001",
		641 => "011001100100001110001",
		642 => "011001100100001110001",
		643 => "011001100100001110001",
		644 => "011001100100001110001",
		645 => "011001100100001110001",
		646 => "011001100100001110001",
		647 => "011001100100001110001",
		648 => "011001100100001110001",
		649 => "011001100100001110001",
		650 => "011001100100001110001",
		651 => "011001100100001110001",
		652 => "011001100100001110001",
		653 => "011001100100001110001",
		654 => "011001100100001110001",
		655 => "011001100100001110001",
		656 => "011001100100001110001",
		657 => "011001100100001110001",
		658 => "011001100100001110001",
		659 => "011001100100001110001",
		660 => "011001100100001110001",
		661 => "011001100100001110001",
		662 => "011001100100001110001",
		663 => "011001100100001110001",
		664 => "011001100100001110001",
		665 => "011001100100001110001",
		666 => "011001100100001110001",
		667 => "011001100100001110001",
		668 => "011001100100001110001",
		669 => "011001100100001110001",
		670 => "011001100100001110001",
		671 => "011001100100001110001",
		672 => "011000101100100010101",
		673 => "011000101100100010101",
		674 => "011000101100100010101",
		675 => "011000101100100010101",
		676 => "011000101100100010101",
		677 => "011000101100100010101",
		678 => "011000101100100010101",
		679 => "011000101100100010101",
		680 => "011000101100100010101",
		681 => "011000101100100010101",
		682 => "011000101100100010101",
		683 => "011000101100100010101",
		684 => "011000101100100010101",
		685 => "011000101100100010101",
		686 => "011000101100100010101",
		687 => "011000101100100010101",
		688 => "011000101100100010101",
		689 => "011000101100100010101",
		690 => "011000101100100010101",
		691 => "011000101100100010101",
		692 => "011000101100100010101",
		693 => "011000101100100010101",
		694 => "011000101100100010101",
		695 => "011000101100100010101",
		696 => "011000101100100010101",
		697 => "011000101100100010101",
		698 => "011000101100100010101",
		699 => "011000101100100010101",
		700 => "011000101100100010101",
		701 => "011000101100100010101",
		702 => "011000101100100010101",
		703 => "011000101100100010101",
		704 => "011000101100100010101",
		705 => "011000101100100010101",
		706 => "011000101100100010101",
		707 => "011000101100100010101",
		708 => "011000101100100010101",
		709 => "011000101100100010101",
		710 => "011000101100100010101",
		711 => "011000101100100010101",
		712 => "011000101100100010101",
		713 => "011000101100100010101",
		714 => "011000101100100010101",
		715 => "011000101100100010101",
		716 => "011000101100100010101",
		717 => "011000101100100010101",
		718 => "011000101100100010101",
		719 => "011000101100100010101",
		720 => "011000101100100010101",
		721 => "011000101100100010101",
		722 => "011000101100100010101",
		723 => "011000101100100010101",
		724 => "011000101100100010101",
		725 => "011000101100100010101",
		726 => "011000101100100010101",
		727 => "011000101100100010101",
		728 => "011000101100100010101",
		729 => "011000101100100010101",
		730 => "011000101100100010101",
		731 => "011000101100100010101",
		732 => "011000101100100010101",
		733 => "011000101100100010101",
		734 => "011000101100100010101",
		735 => "011000101100100010101",
		736 => "011000101100100010101",
		737 => "011000101100100010101",
		738 => "011000101100100010101",
		739 => "011000101100100010101",
		740 => "011000101100100010101",
		741 => "011000101100100010101",
		742 => "011000101100100010101",
		743 => "011000101100100010101",
		744 => "011000101100100010101",
		745 => "011000101100100010101",
		746 => "011000101100100010101",
		747 => "011000101100100010101",
		748 => "011000101100100010101",
		749 => "011000101100100010101",
		750 => "011000101100100010101",
		751 => "011000101100100010101",
		752 => "011000101100100010101",
		753 => "011000101100100010101",
		754 => "011000101100100010101",
		755 => "011000101100100010101",
		756 => "011000101100100010101",
		757 => "011000101100100010101",
		758 => "011000101100100010101",
		759 => "011000101100100010101",
		760 => "011000101100100010101",
		761 => "011000101100100010101",
		762 => "011000101100100010101",
		763 => "011000101100100010101",
		764 => "011000101100100010101",
		765 => "011000101100100010101",
		766 => "011000101100100010101",
		767 => "011000101100100010101",
		768 => "011000101100100110010",
		769 => "011000101100100110010",
		770 => "011000101100100110010",
		771 => "011000101100100110010",
		772 => "011000101100100110010",
		773 => "011000101100100110010",
		774 => "011000101100100110010",
		775 => "011000101100100110010",
		776 => "011000101100100110010",
		777 => "011000101100100110010",
		778 => "011000101100100110010",
		779 => "011000101100100110010",
		780 => "011000101100100110010",
		781 => "011000101100100110010",
		782 => "011000101100100110010",
		783 => "011000101100100110010",
		784 => "011000101100100110010",
		785 => "011000101100100110010",
		786 => "011000101100100110010",
		787 => "011000101100100110010",
		788 => "011000101100100110010",
		789 => "011000101100100110010",
		790 => "011000101100100110010",
		791 => "011000101100100110010",
		792 => "011000101100100110010",
		793 => "011000101100100110010",
		794 => "011000101100100110010",
		795 => "011000101100100110010",
		796 => "011000101100100110010",
		797 => "011000101100100110010",
		798 => "011000101100100110010",
		799 => "011000101100100110010",
		800 => "011000101100100110010",
		801 => "011000101100100110010",
		802 => "011000101100100110010",
		803 => "011000101100100110010",
		804 => "011000101100100110010",
		805 => "011000101100100110010",
		806 => "011000101100100110010",
		807 => "011000101100100110010",
		808 => "011000101100100110010",
		809 => "011000101100100110010",
		810 => "011000101100100110010",
		811 => "011000101100100110010",
		812 => "011000101100100110010",
		813 => "011000101100100110010",
		814 => "011000101100100110010",
		815 => "011000101100100110010",
		816 => "011000101100100110010",
		817 => "011000101100100110010",
		818 => "011000101100100110010",
		819 => "011000101100100110010",
		820 => "011000101100100110010",
		821 => "011000101100100110010",
		822 => "011000101100100110010",
		823 => "011000101100100110010",
		824 => "011000101100100110010",
		825 => "011000101100100110010",
		826 => "011000101100100110010",
		827 => "011000101100100110010",
		828 => "011000101100100110010",
		829 => "011000101100100110010",
		830 => "011000101100100110010",
		831 => "011000101100100110010",
		832 => "011000101100100110010",
		833 => "011000101100100110010",
		834 => "011000101100100110010",
		835 => "011000101100100110010",
		836 => "011000101100100110010",
		837 => "011000101100100110010",
		838 => "011000101100100110010",
		839 => "011000101100100110010",
		840 => "011000101100100110010",
		841 => "011000101100100110010",
		842 => "011000101100100110010",
		843 => "011000101100100110010",
		844 => "011000101100100110010",
		845 => "011000101100100110010",
		846 => "011000101100100110010",
		847 => "011000101100100110010",
		848 => "011000101100100110010",
		849 => "011000101100100110010",
		850 => "011000101100100110010",
		851 => "011000101100100110010",
		852 => "011000101100100110010",
		853 => "011000101100100110010",
		854 => "011000101100100110010",
		855 => "011000101100100110010",
		856 => "011000101100100110010",
		857 => "011000101100100110010",
		858 => "011000101100100110010",
		859 => "011000101100100110010",
		860 => "011000101100100110010",
		861 => "011000101100100110010",
		862 => "011000101100100110010",
		863 => "011000101100100110010");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;