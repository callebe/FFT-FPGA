library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROMFFT1024p_3 is
	Port(
		Adress : in STD_LOGIC;
		reset : in STD_LOGIC;
		Data : out STD_LOGIC_VECTOR (20 downto 0)
		);
end ROMFFT1024p_3;

architecture Behavioral of ROMFFT1024p_3 is

	type ROM is array (863 downto 0) of std_logic_vector(20 downto 0) ;
	-- ROM 4 
	constant ROM_tb : ROM := (
		0 => "001000011110101011000",
		1 => "001000011110101011000",
		2 => "001000011110101011000",
		3 => "011100011110011010000",
		4 => "011100011110011010000",
		5 => "011100011110011010000",
		6 => "011011100100001110111",
		7 => "011011100100001110111",
		8 => "011011100100001110111",
		9 => "011001111100101010000",
		10 => "011001111100101010000",
		11 => "011001111100101010000",
		12 => "001000000100111010010",
		13 => "001000000100111010010",
		14 => "001000000100111010010",
		15 => "011000000101101110010",
		16 => "011000000101101110010",
		17 => "011000000101101110010",
		18 => "011010011101011010000",
		19 => "011010011101011010000",
		20 => "011010011101011010000",
		21 => "011000000100111010011",
		22 => "011000000100111010011",
		23 => "011000000100111010011",
		24 => "011000000100111110001",
		25 => "011000000100111110001",
		26 => "011000000100111110001",
		27 => "011000000100111010110",
		28 => "011000000100111010110",
		29 => "011000000100111010110",
		30 => "011010000100001010010",
		31 => "011010000100001010010",
		32 => "011010000100001010010",
		33 => "001000111100001010011",
		34 => "001000111100001010011",
		35 => "001000111100001010011",
		36 => "011001001100111010000",
		37 => "011001001100111010000",
		38 => "011001001100111010000",
		39 => "011000000100111010000",
		40 => "011000000100111010000",
		41 => "011000000100111010000",
		42 => "011000110100011010011",
		43 => "011000110100011010011",
		44 => "011000110100011010011",
		45 => "001001011100001010011",
		46 => "001001011100001010011",
		47 => "001001011100001010011",
		48 => "011001100100001110000",
		49 => "011001100100001110000",
		50 => "011001100100001110000",
		51 => "011000011100111010000",
		52 => "011000011100111010000",
		53 => "011000011100111010000",
		54 => "001000100100111110001",
		55 => "001000100100111110001",
		56 => "001000100100111110001",
		57 => "001001111100011110010",
		58 => "001001111100011110010",
		59 => "001001111100011110010",
		60 => "011001000100001110001",
		61 => "011001000100001110001",
		62 => "011001000100001110001",
		63 => "011000000100111010001",
		64 => "011000000100111010001",
		65 => "011000000100111010001",
		66 => "011001011100001010100",
		67 => "011001011100001010100",
		68 => "011001011100001010100",
		69 => "011010000100001110001",
		70 => "011010000100001110001",
		71 => "011010000100001110001",
		72 => "011000000101111010010",
		73 => "011000000101111010010",
		74 => "011000000101111010010",
		75 => "011000000101011010100",
		76 => "011000000101011010100",
		77 => "011000000101011010100",
		78 => "011000000101011010101",
		79 => "011000000101011010101",
		80 => "011000000101011010101",
		81 => "011011011101011010000",
		82 => "011011011101011010000",
		83 => "011011011101011010000",
		84 => "011000000101111010011",
		85 => "011000000101111010011",
		86 => "011000000101111010011",
		87 => "011000010101001011000",
		88 => "011000010101001011000",
		89 => "011000010101001011000",
		90 => "011000000110011010110",
		91 => "011000000110011010110",
		92 => "011000000110011010110",
		93 => "011101100100001011011",
		94 => "011101100100001011011",
		95 => "011101100100001011011",
		96 => "011100001110011010000",
		97 => "011100001110011010000",
		98 => "011100001110011010000",
		99 => "001001111100001010111",
		100 => "001001111100001010111",
		101 => "001001111100001010111",
		102 => "001001011100001010110",
		103 => "001001011100001010110",
		104 => "001001011100001010110",
		105 => "011000111100111010000",
		106 => "011000111100111010000",
		107 => "011000111100111010000",
		108 => "001000011100111010001",
		109 => "001000011100111010001",
		110 => "001000011100111010001",
		111 => "011000111100111010000",
		112 => "011000111100111010000",
		113 => "011000111100111010000",
		114 => "011000000100111010000",
		115 => "011000000100111010000",
		116 => "011000000100111010000",
		117 => "011001100100001110000",
		118 => "011001100100001110000",
		119 => "011001100100001110000",
		120 => "011000000100111010010",
		121 => "011000000100111010010",
		122 => "011000000100111010010",
		123 => "011000000101101010011",
		124 => "011000000101101010011",
		125 => "011000000101101010011",
		126 => "011000000101001010001",
		127 => "011000000101001010001",
		128 => "011000000101001010001",
		129 => "111000011101011010011",
		130 => "111000011101011010011",
		131 => "111000011101011010011",
		132 => "001000011100101110011",
		133 => "001000011100101110011",
		134 => "001000011100101110011",
		135 => "011000000101011010111",
		136 => "011000000101011010111",
		137 => "011000000101011010111",
		138 => "011000000101111010011",
		139 => "011000000101111010011",
		140 => "011000000101111010011",
		141 => "011000001100110110110",
		142 => "011000001100110110110",
		143 => "011000001100110110110",
		144 => "001000011110011010111",
		145 => "001000011110011010111",
		146 => "001000011110011010111",
		147 => "011011100100001010011",
		148 => "011011100100001010011",
		149 => "011011100100001010011",
		150 => "011011000100001010010",
		151 => "011011000100001010010",
		152 => "011011000100001010010",
		153 => "011000111100111010000",
		154 => "011000111100111010000",
		155 => "011000111100111010000",
		156 => "011010000100001010100",
		157 => "011010000100001010100",
		158 => "011010000100001010100",
		159 => "011000111100111010000",
		160 => "011000111100111010000",
		161 => "011000111100111010000",
		162 => "011001100100001110000",
		163 => "011001100100001110000",
		164 => "011001100100001110000",
		165 => "001000011100111010000",
		166 => "001000011100111010000",
		167 => "001000011100111010000",
		168 => "011000000101101010001",
		169 => "011000000101101010001",
		170 => "011000000101101010001",
		171 => "011000000101101010011",
		172 => "011000000101101010011",
		173 => "011000000101101010011",
		174 => "011000000101001010001",
		175 => "011000000101001010001",
		176 => "011000000101001010001",
		177 => "011000001101010010011",
		178 => "011000001101010010011",
		179 => "011000001101010010011",
		180 => "011001100100011010000",
		181 => "011001100100011010000",
		182 => "011001100100011010000",
		183 => "011000010100101011000",
		184 => "011000010100101011000",
		185 => "011000010100101011000",
		186 => "001001111101111010000",
		187 => "001001111101111010000",
		188 => "001001111101111010000",
		189 => "011000001100110110110",
		190 => "011000001100110110110",
		191 => "011000001100110110110",
		192 => "011011101110001010000",
		193 => "011011101110001010000",
		194 => "011011101110001010000",
		195 => "001001100101101110000",
		196 => "001001100101101110000",
		197 => "001001100101101110000",
		198 => "011000001101100010011",
		199 => "011000001101100010011",
		200 => "011000001101100010011",
		201 => "011000001100101010110",
		202 => "011000001100101010110",
		203 => "011000001100101010110",
		204 => "011000101100101010100",
		205 => "011000101100101010100",
		206 => "011000101100101010100",
		207 => "011000000100111010001",
		208 => "011000000100111010001",
		209 => "011000000100111010001",
		210 => "011000000101011010010",
		211 => "011000000101011010010",
		212 => "011000000101011010010",
		213 => "001001111110001010000",
		214 => "001001111110001010000",
		215 => "001001111110001010000",
		216 => "001000011110001010110",
		217 => "001000011110001010110",
		218 => "001000011110001010110",
		219 => "001000010100111010110",
		220 => "001000010100111010110",
		221 => "001000010100111010110",
		222 => "011000001101100010011",
		223 => "011000001101100010011",
		224 => "011000001101100010011",
		225 => "001000111100011110011",
		226 => "001000111100011110011",
		227 => "001000111100011110011",
		228 => "011001000100001110100",
		229 => "011001000100001110100",
		230 => "011001000100001110100",
		231 => "011000000100111010001",
		232 => "011000000100111010001",
		233 => "011000000100111010001",
		234 => "011000000101011010010",
		235 => "011000000101011010010",
		236 => "011000000101011010010",
		237 => "001001111110001010000",
		238 => "001001111110001010000",
		239 => "001001111110001010000",
		240 => "011011101110001010000",
		241 => "011011101110001010000",
		242 => "011011101110001010000",
		243 => "001001100101101110000",
		244 => "001001100101101110000",
		245 => "001001100101101110000",
		246 => "011000001101100010011",
		247 => "011000001101100010011",
		248 => "011000001101100010011",
		249 => "011000001100101010110",
		250 => "011000001100101010110",
		251 => "011000001100101010110",
		252 => "011000101100101010100",
		253 => "011000101100101010100",
		254 => "011000101100101010100",
		255 => "011000000100111010001",
		256 => "011000000100111010001",
		257 => "011000000100111010001",
		258 => "011000000101011010010",
		259 => "011000000101011010010",
		260 => "011000000101011010010",
		261 => "001001111110001010000",
		262 => "001001111110001010000",
		263 => "001001111110001010000",
		264 => "001000011110001010110",
		265 => "001000011110001010110",
		266 => "001000011110001010110",
		267 => "001000010100111010110",
		268 => "001000010100111010110",
		269 => "001000010100111010110",
		270 => "011000001101100010011",
		271 => "011000001101100010011",
		272 => "011000001101100010011",
		273 => "001000111100011110011",
		274 => "001000111100011110011",
		275 => "001000111100011110011",
		276 => "011001000100001110100",
		277 => "011001000100001110100",
		278 => "011001000100001110100",
		279 => "011000000100111010001",
		280 => "011000000100111010001",
		281 => "011000000100111010001",
		282 => "011000000101011010010",
		283 => "011000000101011010010",
		284 => "011000000101011010010",
		285 => "001001111110001010000",
		286 => "001001111110001010000",
		287 => "001001111110001010000",
		288 => "011000000101110011001",
		289 => "011000000101110011001",
		290 => "011000000101110011001",
		291 => "001011011100001010111",
		292 => "001011011100001010111",
		293 => "001011011100001010111",
		294 => "011000000101101010011",
		295 => "011000000101101010011",
		296 => "011000000101101010011",
		297 => "011000001110100010101",
		298 => "011000001110100010101",
		299 => "011000001110100010101",
		300 => "011000000101110011001",
		301 => "011000000101110011001",
		302 => "011000000101110011001",
		303 => "011000111100111010000",
		304 => "011000111100111010000",
		305 => "011000111100111010000",
		306 => "011000000101101010011",
		307 => "011000000101101010011",
		308 => "011000000101101010011",
		309 => "011000001110100010101",
		310 => "011000001110100010101",
		311 => "011000001110100010101",
		312 => "011000000101110011001",
		313 => "011000000101110011001",
		314 => "011000000101110011001",
		315 => "001011011100001010111",
		316 => "001011011100001010111",
		317 => "001011011100001010111",
		318 => "011000000101101010011",
		319 => "011000000101101010011",
		320 => "011000000101101010011",
		321 => "011000001110100010101",
		322 => "011000001110100010101",
		323 => "011000001110100010101",
		324 => "011000000101110011001",
		325 => "011000000101110011001",
		326 => "011000000101110011001",
		327 => "011000111100111010000",
		328 => "011000111100111010000",
		329 => "011000111100111010000",
		330 => "011000000101101010011",
		331 => "011000000101101010011",
		332 => "011000000101101010011",
		333 => "011000001110100010101",
		334 => "011000001110100010101",
		335 => "011000001110100010101",
		336 => "011000000101110011001",
		337 => "011000000101110011001",
		338 => "011000000101110011001",
		339 => "001011011100001010111",
		340 => "001011011100001010111",
		341 => "001011011100001010111",
		342 => "011000000101101010011",
		343 => "011000000101101010011",
		344 => "011000000101101010011",
		345 => "011000001110100010101",
		346 => "011000001110100010101",
		347 => "011000001110100010101",
		348 => "011000000101110011001",
		349 => "011000000101110011001",
		350 => "011000000101110011001",
		351 => "011000111100111010000",
		352 => "011000111100111010000",
		353 => "011000111100111010000",
		354 => "011000000101101010011",
		355 => "011000000101101010011",
		356 => "011000000101101010011",
		357 => "011000001110100010101",
		358 => "011000001110100010101",
		359 => "011000001110100010101",
		360 => "011000000101110011001",
		361 => "011000000101110011001",
		362 => "011000000101110011001",
		363 => "001011011100001010111",
		364 => "001011011100001010111",
		365 => "001011011100001010111",
		366 => "011000000101101010011",
		367 => "011000000101101010011",
		368 => "011000000101101010011",
		369 => "011000001110100010101",
		370 => "011000001110100010101",
		371 => "011000001110100010101",
		372 => "011000000101110011001",
		373 => "011000000101110011001",
		374 => "011000000101110011001",
		375 => "011000111100111010000",
		376 => "011000111100111010000",
		377 => "011000111100111010000",
		378 => "011000000101101010011",
		379 => "011000000101101010011",
		380 => "011000000101101010011",
		381 => "011000001110100010101",
		382 => "011000001110100010101",
		383 => "011000001110100010101",
		384 => "001010111100001010101",
		385 => "001010111100001010101",
		386 => "001010111100001010101",
		387 => "011001011100001010100",
		388 => "011001011100001010100",
		389 => "011001011100001010100",
		390 => "011010100100001010101",
		391 => "011010100100001010101",
		392 => "011010100100001010101",
		393 => "011010000100001110010",
		394 => "011010000100001110010",
		395 => "011010000100001110010",
		396 => "001010111100001010101",
		397 => "001010111100001010101",
		398 => "001010111100001010101",
		399 => "011001011100001010100",
		400 => "011001011100001010100",
		401 => "011001011100001010100",
		402 => "011010100100001010101",
		403 => "011010100100001010101",
		404 => "011010100100001010101",
		405 => "011010000100001110010",
		406 => "011010000100001110010",
		407 => "011010000100001110010",
		408 => "001010111100001010101",
		409 => "001010111100001010101",
		410 => "001010111100001010101",
		411 => "011001011100001010100",
		412 => "011001011100001010100",
		413 => "011001011100001010100",
		414 => "011010100100001010101",
		415 => "011010100100001010101",
		416 => "011010100100001010101",
		417 => "011010000100001110010",
		418 => "011010000100001110010",
		419 => "011010000100001110010",
		420 => "001010111100001010101",
		421 => "001010111100001010101",
		422 => "001010111100001010101",
		423 => "011001011100001010100",
		424 => "011001011100001010100",
		425 => "011001011100001010100",
		426 => "011010100100001010101",
		427 => "011010100100001010101",
		428 => "011010100100001010101",
		429 => "011010000100001110010",
		430 => "011010000100001110010",
		431 => "011010000100001110010",
		432 => "001010111100001010101",
		433 => "001010111100001010101",
		434 => "001010111100001010101",
		435 => "011001011100001010100",
		436 => "011001011100001010100",
		437 => "011001011100001010100",
		438 => "011010100100001010101",
		439 => "011010100100001010101",
		440 => "011010100100001010101",
		441 => "011010000100001110010",
		442 => "011010000100001110010",
		443 => "011010000100001110010",
		444 => "001010111100001010101",
		445 => "001010111100001010101",
		446 => "001010111100001010101",
		447 => "011001011100001010100",
		448 => "011001011100001010100",
		449 => "011001011100001010100",
		450 => "011010100100001010101",
		451 => "011010100100001010101",
		452 => "011010100100001010101",
		453 => "011010000100001110010",
		454 => "011010000100001110010",
		455 => "011010000100001110010",
		456 => "001010111100001010101",
		457 => "001010111100001010101",
		458 => "001010111100001010101",
		459 => "011001011100001010100",
		460 => "011001011100001010100",
		461 => "011001011100001010100",
		462 => "011010100100001010101",
		463 => "011010100100001010101",
		464 => "011010100100001010101",
		465 => "011010000100001110010",
		466 => "011010000100001110010",
		467 => "011010000100001110010",
		468 => "001010111100001010101",
		469 => "001010111100001010101",
		470 => "001010111100001010101",
		471 => "011001011100001010100",
		472 => "011001011100001010100",
		473 => "011001011100001010100",
		474 => "011010100100001010101",
		475 => "011010100100001010101",
		476 => "011010100100001010101",
		477 => "011010000100001110010",
		478 => "011010000100001110010",
		479 => "011010000100001110010",
		480 => "011000001101100010011",
		481 => "011000001101100010011",
		482 => "011000001101100010011",
		483 => "011000001101100010011",
		484 => "011000001101100010011",
		485 => "011000001101100010011",
		486 => "011000001101100010011",
		487 => "011000001101100010011",
		488 => "011000001101100010011",
		489 => "011000001101100010011",
		490 => "011000001101100010011",
		491 => "011000001101100010011",
		492 => "011000001101100010011",
		493 => "011000001101100010011",
		494 => "011000001101100010011",
		495 => "011000001101100010011",
		496 => "011000001101100010011",
		497 => "011000001101100010011",
		498 => "011000001101100010011",
		499 => "011000001101100010011",
		500 => "011000001101100010011",
		501 => "011000001101100010011",
		502 => "011000001101100010011",
		503 => "011000001101100010011",
		504 => "011000001101100010011",
		505 => "011000001101100010011",
		506 => "011000001101100010011",
		507 => "011000001101100010011",
		508 => "011000001101100010011",
		509 => "011000001101100010011",
		510 => "011000001101100010011",
		511 => "011000001101100010011",
		512 => "011000001101100010011",
		513 => "011000001101100010011",
		514 => "011000001101100010011",
		515 => "011000001101100010011",
		516 => "011000001101100010011",
		517 => "011000001101100010011",
		518 => "011000001101100010011",
		519 => "011000001101100010011",
		520 => "011000001101100010011",
		521 => "011000001101100010011",
		522 => "011000001101100010011",
		523 => "011000001101100010011",
		524 => "011000001101100010011",
		525 => "011000001101100010011",
		526 => "011000001101100010011",
		527 => "011000001101100010011",
		528 => "011000001101100010011",
		529 => "011000001101100010011",
		530 => "011000001101100010011",
		531 => "011000001101100010011",
		532 => "011000001101100010011",
		533 => "011000001101100010011",
		534 => "011000001101100010011",
		535 => "011000001101100010011",
		536 => "011000001101100010011",
		537 => "011000001101100010011",
		538 => "011000001101100010011",
		539 => "011000001101100010011",
		540 => "011000001101100010011",
		541 => "011000001101100010011",
		542 => "011000001101100010011",
		543 => "011000001101100010011",
		544 => "011000001101100010011",
		545 => "011000001101100010011",
		546 => "011000001101100010011",
		547 => "011000001101100010011",
		548 => "011000001101100010011",
		549 => "011000001101100010011",
		550 => "011000001101100010011",
		551 => "011000001101100010011",
		552 => "011000001101100010011",
		553 => "011000001101100010011",
		554 => "011000001101100010011",
		555 => "011000001101100010011",
		556 => "011000001101100010011",
		557 => "011000001101100010011",
		558 => "011000001101100010011",
		559 => "011000001101100010011",
		560 => "011000001101100010011",
		561 => "011000001101100010011",
		562 => "011000001101100010011",
		563 => "011000001101100010011",
		564 => "011000001101100010011",
		565 => "011000001101100010011",
		566 => "011000001101100010011",
		567 => "011000001101100010011",
		568 => "011000001101100010011",
		569 => "011000001101100010011",
		570 => "011000001101100010011",
		571 => "011000001101100010011",
		572 => "011000001101100010011",
		573 => "011000001101100010011",
		574 => "011000001101100010011",
		575 => "011000001101100010011",
		576 => "011001100100001110001",
		577 => "011001100100001110001",
		578 => "011001100100001110001",
		579 => "011001100100001110001",
		580 => "011001100100001110001",
		581 => "011001100100001110001",
		582 => "011001100100001110001",
		583 => "011001100100001110001",
		584 => "011001100100001110001",
		585 => "011001100100001110001",
		586 => "011001100100001110001",
		587 => "011001100100001110001",
		588 => "011001100100001110001",
		589 => "011001100100001110001",
		590 => "011001100100001110001",
		591 => "011001100100001110001",
		592 => "011001100100001110001",
		593 => "011001100100001110001",
		594 => "011001100100001110001",
		595 => "011001100100001110001",
		596 => "011001100100001110001",
		597 => "011001100100001110001",
		598 => "011001100100001110001",
		599 => "011001100100001110001",
		600 => "011001100100001110001",
		601 => "011001100100001110001",
		602 => "011001100100001110001",
		603 => "011001100100001110001",
		604 => "011001100100001110001",
		605 => "011001100100001110001",
		606 => "011001100100001110001",
		607 => "011001100100001110001",
		608 => "011001100100001110001",
		609 => "011001100100001110001",
		610 => "011001100100001110001",
		611 => "011001100100001110001",
		612 => "011001100100001110001",
		613 => "011001100100001110001",
		614 => "011001100100001110001",
		615 => "011001100100001110001",
		616 => "011001100100001110001",
		617 => "011001100100001110001",
		618 => "011001100100001110001",
		619 => "011001100100001110001",
		620 => "011001100100001110001",
		621 => "011001100100001110001",
		622 => "011001100100001110001",
		623 => "011001100100001110001",
		624 => "011001100100001110001",
		625 => "011001100100001110001",
		626 => "011001100100001110001",
		627 => "011001100100001110001",
		628 => "011001100100001110001",
		629 => "011001100100001110001",
		630 => "011001100100001110001",
		631 => "011001100100001110001",
		632 => "011001100100001110001",
		633 => "011001100100001110001",
		634 => "011001100100001110001",
		635 => "011001100100001110001",
		636 => "011001100100001110001",
		637 => "011001100100001110001",
		638 => "011001100100001110001",
		639 => "011001100100001110001",
		640 => "011001100100001110001",
		641 => "011001100100001110001",
		642 => "011001100100001110001",
		643 => "011001100100001110001",
		644 => "011001100100001110001",
		645 => "011001100100001110001",
		646 => "011001100100001110001",
		647 => "011001100100001110001",
		648 => "011001100100001110001",
		649 => "011001100100001110001",
		650 => "011001100100001110001",
		651 => "011001100100001110001",
		652 => "011001100100001110001",
		653 => "011001100100001110001",
		654 => "011001100100001110001",
		655 => "011001100100001110001",
		656 => "011001100100001110001",
		657 => "011001100100001110001",
		658 => "011001100100001110001",
		659 => "011001100100001110001",
		660 => "011001100100001110001",
		661 => "011001100100001110001",
		662 => "011001100100001110001",
		663 => "011001100100001110001",
		664 => "011001100100001110001",
		665 => "011001100100001110001",
		666 => "011001100100001110001",
		667 => "011001100100001110001",
		668 => "011001100100001110001",
		669 => "011001100100001110001",
		670 => "011001100100001110001",
		671 => "011001100100001110001",
		672 => "011000101100100010101",
		673 => "011000101100100010101",
		674 => "011000101100100010101",
		675 => "011000101100100010101",
		676 => "011000101100100010101",
		677 => "011000101100100010101",
		678 => "011000101100100010101",
		679 => "011000101100100010101",
		680 => "011000101100100010101",
		681 => "011000101100100010101",
		682 => "011000101100100010101",
		683 => "011000101100100010101",
		684 => "011000101100100010101",
		685 => "011000101100100010101",
		686 => "011000101100100010101",
		687 => "011000101100100010101",
		688 => "011000101100100010101",
		689 => "011000101100100010101",
		690 => "011000101100100010101",
		691 => "011000101100100010101",
		692 => "011000101100100010101",
		693 => "011000101100100010101",
		694 => "011000101100100010101",
		695 => "011000101100100010101",
		696 => "011000101100100010101",
		697 => "011000101100100010101",
		698 => "011000101100100010101",
		699 => "011000101100100010101",
		700 => "011000101100100010101",
		701 => "011000101100100010101",
		702 => "011000101100100010101",
		703 => "011000101100100010101",
		704 => "011000101100100010101",
		705 => "011000101100100010101",
		706 => "011000101100100010101",
		707 => "011000101100100010101",
		708 => "011000101100100010101",
		709 => "011000101100100010101",
		710 => "011000101100100010101",
		711 => "011000101100100010101",
		712 => "011000101100100010101",
		713 => "011000101100100010101",
		714 => "011000101100100010101",
		715 => "011000101100100010101",
		716 => "011000101100100010101",
		717 => "011000101100100010101",
		718 => "011000101100100010101",
		719 => "011000101100100010101",
		720 => "011000101100100010101",
		721 => "011000101100100010101",
		722 => "011000101100100010101",
		723 => "011000101100100010101",
		724 => "011000101100100010101",
		725 => "011000101100100010101",
		726 => "011000101100100010101",
		727 => "011000101100100010101",
		728 => "011000101100100010101",
		729 => "011000101100100010101",
		730 => "011000101100100010101",
		731 => "011000101100100010101",
		732 => "011000101100100010101",
		733 => "011000101100100010101",
		734 => "011000101100100010101",
		735 => "011000101100100010101",
		736 => "011000101100100010101",
		737 => "011000101100100010101",
		738 => "011000101100100010101",
		739 => "011000101100100010101",
		740 => "011000101100100010101",
		741 => "011000101100100010101",
		742 => "011000101100100010101",
		743 => "011000101100100010101",
		744 => "011000101100100010101",
		745 => "011000101100100010101",
		746 => "011000101100100010101",
		747 => "011000101100100010101",
		748 => "011000101100100010101",
		749 => "011000101100100010101",
		750 => "011000101100100010101",
		751 => "011000101100100010101",
		752 => "011000101100100010101",
		753 => "011000101100100010101",
		754 => "011000101100100010101",
		755 => "011000101100100010101",
		756 => "011000101100100010101",
		757 => "011000101100100010101",
		758 => "011000101100100010101",
		759 => "011000101100100010101",
		760 => "011000101100100010101",
		761 => "011000101100100010101",
		762 => "011000101100100010101",
		763 => "011000101100100010101",
		764 => "011000101100100010101",
		765 => "011000101100100010101",
		766 => "011000101100100010101",
		767 => "011000101100100010101",
		768 => "011000101100100110010",
		769 => "011000101100100110010",
		770 => "011000101100100110010",
		771 => "011000101100100110010",
		772 => "011000101100100110010",
		773 => "011000101100100110010",
		774 => "011000101100100110010",
		775 => "011000101100100110010",
		776 => "011000101100100110010",
		777 => "011000101100100110010",
		778 => "011000101100100110010",
		779 => "011000101100100110010",
		780 => "011000101100100110010",
		781 => "011000101100100110010",
		782 => "011000101100100110010",
		783 => "011000101100100110010",
		784 => "011000101100100110010",
		785 => "011000101100100110010",
		786 => "011000101100100110010",
		787 => "011000101100100110010",
		788 => "011000101100100110010",
		789 => "011000101100100110010",
		790 => "011000101100100110010",
		791 => "011000101100100110010",
		792 => "011000101100100110010",
		793 => "011000101100100110010",
		794 => "011000101100100110010",
		795 => "011000101100100110010",
		796 => "011000101100100110010",
		797 => "011000101100100110010",
		798 => "011000101100100110010",
		799 => "011000101100100110010",
		800 => "011000101100100110010",
		801 => "011000101100100110010",
		802 => "011000101100100110010",
		803 => "011000101100100110010",
		804 => "011000101100100110010",
		805 => "011000101100100110010",
		806 => "011000101100100110010",
		807 => "011000101100100110010",
		808 => "011000101100100110010",
		809 => "011000101100100110010",
		810 => "011000101100100110010",
		811 => "011000101100100110010",
		812 => "011000101100100110010",
		813 => "011000101100100110010",
		814 => "011000101100100110010",
		815 => "011000101100100110010",
		816 => "011000101100100110010",
		817 => "011000101100100110010",
		818 => "011000101100100110010",
		819 => "011000101100100110010",
		820 => "011000101100100110010",
		821 => "011000101100100110010",
		822 => "011000101100100110010",
		823 => "011000101100100110010",
		824 => "011000101100100110010",
		825 => "011000101100100110010",
		826 => "011000101100100110010",
		827 => "011000101100100110010",
		828 => "011000101100100110010",
		829 => "011000101100100110010",
		830 => "011000101100100110010",
		831 => "011000101100100110010",
		832 => "011000101100100110010",
		833 => "011000101100100110010",
		834 => "011000101100100110010",
		835 => "011000101100100110010",
		836 => "011000101100100110010",
		837 => "011000101100100110010",
		838 => "011000101100100110010",
		839 => "011000101100100110010",
		840 => "011000101100100110010",
		841 => "011000101100100110010",
		842 => "011000101100100110010",
		843 => "011000101100100110010",
		844 => "011000101100100110010",
		845 => "011000101100100110010",
		846 => "011000101100100110010",
		847 => "011000101100100110010",
		848 => "011000101100100110010",
		849 => "011000101100100110010",
		850 => "011000101100100110010",
		851 => "011000101100100110010",
		852 => "011000101100100110010",
		853 => "011000101100100110010",
		854 => "011000101100100110010",
		855 => "011000101100100110010",
		856 => "011000101100100110010",
		857 => "011000101100100110010",
		858 => "011000101100100110010",
		859 => "011000101100100110010",
		860 => "011000101100100110010",
		861 => "011000101100100110010",
		862 => "011000101100100110010",
		863 => "011000101100100110010");

	begin
		--Process to acess Data
		process(Adress, reset)

			variable Counter : integer range 510 downto 0 := 0;

		begin

		Data <= Rom_tb(Counter);
		if(reset = '1')then
			Counter := 0;

		elsif(Adress'event and Adress = '1') then
			Counter := Counter + 1;

		end if;

	end process;

end Behavioral;